/////////////////////////////////////////////////////////////////////////////////
// Company       : �人о·��Ƽ����޹�˾
//                 http://xiaomeige.taobao.com
// Web           : http://www.corecourse.cn
// 
// Create Date   : 2019/05/01 00:00:00
// Module Name   : rom_image
// Description   : ͼ��romģ��
// 
// Dependencies  : 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
/////////////////////////////////////////////////////////////////////////////////

module rom_image(
  input             clk ,
  input      [15:0] addr,
  output reg [15:0] dout
);

reg [15:0] rom [65535:0];

initial begin
  rom[00000] = 16'hffff;
  rom[00001] = 16'hffff;
  rom[00002] = 16'hffff;
  rom[00003] = 16'hffff;
  rom[00004] = 16'hffff;
  rom[00005] = 16'hffff;
  rom[00006] = 16'hffff;
  rom[00007] = 16'hffff;
  rom[00008] = 16'hffff;
  rom[00009] = 16'hffff;
  rom[00010] = 16'hffff;
  rom[00011] = 16'hffff;
  rom[00012] = 16'hffff;
  rom[00013] = 16'hffff;
  rom[00014] = 16'hffff;
  rom[00015] = 16'hffff;
  rom[00016] = 16'hffff;
  rom[00017] = 16'hffff;
  rom[00018] = 16'hffff;
  rom[00019] = 16'hffff;
  rom[00020] = 16'hffff;
  rom[00021] = 16'hffff;
  rom[00022] = 16'hffff;
  rom[00023] = 16'hffff;
  rom[00024] = 16'hffff;
  rom[00025] = 16'hffff;
  rom[00026] = 16'hffff;
  rom[00027] = 16'hffff;
  rom[00028] = 16'hffff;
  rom[00029] = 16'hffff;
  rom[00030] = 16'hffff;
  rom[00031] = 16'hffff;
  rom[00032] = 16'hffff;
  rom[00033] = 16'hffff;
  rom[00034] = 16'hffff;
  rom[00035] = 16'hffff;
  rom[00036] = 16'hffff;
  rom[00037] = 16'hffff;
  rom[00038] = 16'hffff;
  rom[00039] = 16'hffff;
  rom[00040] = 16'hffff;
  rom[00041] = 16'hffff;
  rom[00042] = 16'hffff;
  rom[00043] = 16'hffff;
  rom[00044] = 16'hffff;
  rom[00045] = 16'hffff;
  rom[00046] = 16'hffff;
  rom[00047] = 16'hffff;
  rom[00048] = 16'hffff;
  rom[00049] = 16'hffff;
  rom[00050] = 16'hffff;
  rom[00051] = 16'hffff;
  rom[00052] = 16'hffff;
  rom[00053] = 16'hffff;
  rom[00054] = 16'hffff;
  rom[00055] = 16'hffff;
  rom[00056] = 16'hffff;
  rom[00057] = 16'hffff;
  rom[00058] = 16'hffff;
  rom[00059] = 16'hffff;
  rom[00060] = 16'hffff;
  rom[00061] = 16'hffff;
  rom[00062] = 16'hffff;
  rom[00063] = 16'hffff;
  rom[00064] = 16'hffdf;
  rom[00065] = 16'hffff;
  rom[00066] = 16'hffff;
  rom[00067] = 16'hffff;
  rom[00068] = 16'hffff;
  rom[00069] = 16'hffff;
  rom[00070] = 16'hffff;
  rom[00071] = 16'hffff;
  rom[00072] = 16'hffff;
  rom[00073] = 16'hffff;
  rom[00074] = 16'hffff;
  rom[00075] = 16'hffff;
  rom[00076] = 16'hffff;
  rom[00077] = 16'hffff;
  rom[00078] = 16'hffff;
  rom[00079] = 16'hffff;
  rom[00080] = 16'hffff;
  rom[00081] = 16'hffff;
  rom[00082] = 16'hffff;
  rom[00083] = 16'hffff;
  rom[00084] = 16'hffdf;
  rom[00085] = 16'hffff;
  rom[00086] = 16'hffde;
  rom[00087] = 16'hffff;
  rom[00088] = 16'hffbd;
  rom[00089] = 16'hde78;
  rom[00090] = 16'hc593;
  rom[00091] = 16'hcd72;
  rom[00092] = 16'hc552;
  rom[00093] = 16'hf6d8;
  rom[00094] = 16'hf719;
  rom[00095] = 16'h6288;
  rom[00096] = 16'h1880;
  rom[00097] = 16'h18c1;
  rom[00098] = 16'h2143;
  rom[00099] = 16'had95;
  rom[00100] = 16'hf7ff;
  rom[00101] = 16'hffff;
  rom[00102] = 16'hffbf;
  rom[00103] = 16'hffff;
  rom[00104] = 16'hffdf;
  rom[00105] = 16'hffff;
  rom[00106] = 16'hffdf;
  rom[00107] = 16'hffff;
  rom[00108] = 16'hffdf;
  rom[00109] = 16'hffff;
  rom[00110] = 16'hfffe;
  rom[00111] = 16'hffff;
  rom[00112] = 16'hffff;
  rom[00113] = 16'hffff;
  rom[00114] = 16'hffff;
  rom[00115] = 16'hffff;
  rom[00116] = 16'hffff;
  rom[00117] = 16'hffff;
  rom[00118] = 16'hffff;
  rom[00119] = 16'hffff;
  rom[00120] = 16'hffff;
  rom[00121] = 16'hffff;
  rom[00122] = 16'hffff;
  rom[00123] = 16'hffff;
  rom[00124] = 16'hffff;
  rom[00125] = 16'hffff;
  rom[00126] = 16'hffff;
  rom[00127] = 16'hffff;
  rom[00128] = 16'hffff;
  rom[00129] = 16'hffff;
  rom[00130] = 16'hffff;
  rom[00131] = 16'hffff;
  rom[00132] = 16'hffff;
  rom[00133] = 16'hffff;
  rom[00134] = 16'hffdf;
  rom[00135] = 16'hffff;
  rom[00136] = 16'hf7be;
  rom[00137] = 16'hffff;
  rom[00138] = 16'hffdf;
  rom[00139] = 16'hffff;
  rom[00140] = 16'hffff;
  rom[00141] = 16'hffff;
  rom[00142] = 16'hffff;
  rom[00143] = 16'hffff;
  rom[00144] = 16'hffff;
  rom[00145] = 16'hffff;
  rom[00146] = 16'hffff;
  rom[00147] = 16'hffff;
  rom[00148] = 16'hffff;
  rom[00149] = 16'hffff;
  rom[00150] = 16'hffff;
  rom[00151] = 16'hffff;
  rom[00152] = 16'hffff;
  rom[00153] = 16'hffff;
  rom[00154] = 16'hffff;
  rom[00155] = 16'hffff;
  rom[00156] = 16'hffff;
  rom[00157] = 16'hffff;
  rom[00158] = 16'hffff;
  rom[00159] = 16'hffff;
  rom[00160] = 16'hffff;
  rom[00161] = 16'hffff;
  rom[00162] = 16'hffff;
  rom[00163] = 16'hffff;
  rom[00164] = 16'hffff;
  rom[00165] = 16'hffff;
  rom[00166] = 16'hffff;
  rom[00167] = 16'hffff;
  rom[00168] = 16'hffff;
  rom[00169] = 16'hffff;
  rom[00170] = 16'hffff;
  rom[00171] = 16'hffff;
  rom[00172] = 16'hffff;
  rom[00173] = 16'hffff;
  rom[00174] = 16'hffff;
  rom[00175] = 16'hffff;
  rom[00176] = 16'hffff;
  rom[00177] = 16'hffff;
  rom[00178] = 16'hffff;
  rom[00179] = 16'hffff;
  rom[00180] = 16'hffff;
  rom[00181] = 16'hffff;
  rom[00182] = 16'hffff;
  rom[00183] = 16'hffff;
  rom[00184] = 16'hffff;
  rom[00185] = 16'hffff;
  rom[00186] = 16'hffff;
  rom[00187] = 16'hffff;
  rom[00188] = 16'hffff;
  rom[00189] = 16'hffff;
  rom[00190] = 16'hffff;
  rom[00191] = 16'hffff;
  rom[00192] = 16'hffff;
  rom[00193] = 16'hffff;
  rom[00194] = 16'hffff;
  rom[00195] = 16'hffff;
  rom[00196] = 16'hffff;
  rom[00197] = 16'hffff;
  rom[00198] = 16'hffff;
  rom[00199] = 16'hffff;
  rom[00200] = 16'hffff;
  rom[00201] = 16'hffff;
  rom[00202] = 16'hffff;
  rom[00203] = 16'hffff;
  rom[00204] = 16'hffff;
  rom[00205] = 16'hffff;
  rom[00206] = 16'hffff;
  rom[00207] = 16'hffff;
  rom[00208] = 16'hffff;
  rom[00209] = 16'hffff;
  rom[00210] = 16'hffff;
  rom[00211] = 16'hffff;
  rom[00212] = 16'hffff;
  rom[00213] = 16'hffff;
  rom[00214] = 16'hffff;
  rom[00215] = 16'hffff;
  rom[00216] = 16'hffff;
  rom[00217] = 16'hffff;
  rom[00218] = 16'hffff;
  rom[00219] = 16'hffff;
  rom[00220] = 16'hffff;
  rom[00221] = 16'hffff;
  rom[00222] = 16'hffff;
  rom[00223] = 16'hffff;
  rom[00224] = 16'hffff;
  rom[00225] = 16'hffff;
  rom[00226] = 16'hffff;
  rom[00227] = 16'hffff;
  rom[00228] = 16'hffff;
  rom[00229] = 16'hffff;
  rom[00230] = 16'hffff;
  rom[00231] = 16'hffff;
  rom[00232] = 16'hffff;
  rom[00233] = 16'hffff;
  rom[00234] = 16'hffff;
  rom[00235] = 16'hffff;
  rom[00236] = 16'hffff;
  rom[00237] = 16'hffff;
  rom[00238] = 16'hffff;
  rom[00239] = 16'hffff;
  rom[00240] = 16'hffff;
  rom[00241] = 16'hffff;
  rom[00242] = 16'hffff;
  rom[00243] = 16'hffff;
  rom[00244] = 16'hffff;
  rom[00245] = 16'hffff;
  rom[00246] = 16'hffff;
  rom[00247] = 16'hffff;
  rom[00248] = 16'hffff;
  rom[00249] = 16'hffff;
  rom[00250] = 16'hffff;
  rom[00251] = 16'hffff;
  rom[00252] = 16'hffff;
  rom[00253] = 16'hffff;
  rom[00254] = 16'hffff;
  rom[00255] = 16'hffff;
  rom[00256] = 16'hffff;
  rom[00257] = 16'hffff;
  rom[00258] = 16'hffff;
  rom[00259] = 16'hffff;
  rom[00260] = 16'hffff;
  rom[00261] = 16'hffff;
  rom[00262] = 16'hffff;
  rom[00263] = 16'hffff;
  rom[00264] = 16'hffff;
  rom[00265] = 16'hffff;
  rom[00266] = 16'hffff;
  rom[00267] = 16'hffff;
  rom[00268] = 16'hffff;
  rom[00269] = 16'hffff;
  rom[00270] = 16'hffff;
  rom[00271] = 16'hffff;
  rom[00272] = 16'hffff;
  rom[00273] = 16'hffff;
  rom[00274] = 16'hffff;
  rom[00275] = 16'hffff;
  rom[00276] = 16'hffff;
  rom[00277] = 16'hffff;
  rom[00278] = 16'hffff;
  rom[00279] = 16'hffff;
  rom[00280] = 16'hffff;
  rom[00281] = 16'hffff;
  rom[00282] = 16'hffff;
  rom[00283] = 16'hffff;
  rom[00284] = 16'hffff;
  rom[00285] = 16'hffff;
  rom[00286] = 16'hffff;
  rom[00287] = 16'hffde;
  rom[00288] = 16'hffff;
  rom[00289] = 16'h946f;
  rom[00290] = 16'h8b8a;
  rom[00291] = 16'h9baa;
  rom[00292] = 16'h9baa;
  rom[00293] = 16'h7265;
  rom[00294] = 16'h82e7;
  rom[00295] = 16'h30e1;
  rom[00296] = 16'h3101;
  rom[00297] = 16'h18c0;
  rom[00298] = 16'h20e2;
  rom[00299] = 16'h7bef;
  rom[00300] = 16'hffff;
  rom[00301] = 16'hffff;
  rom[00302] = 16'hffff;
  rom[00303] = 16'hffff;
  rom[00304] = 16'hffff;
  rom[00305] = 16'hffff;
  rom[00306] = 16'hffff;
  rom[00307] = 16'hffff;
  rom[00308] = 16'hffff;
  rom[00309] = 16'hffff;
  rom[00310] = 16'hffff;
  rom[00311] = 16'hffff;
  rom[00312] = 16'hffff;
  rom[00313] = 16'hffff;
  rom[00314] = 16'hffff;
  rom[00315] = 16'hffff;
  rom[00316] = 16'hffff;
  rom[00317] = 16'hffff;
  rom[00318] = 16'hffff;
  rom[00319] = 16'hffff;
  rom[00320] = 16'hffff;
  rom[00321] = 16'hffff;
  rom[00322] = 16'hffff;
  rom[00323] = 16'hffff;
  rom[00324] = 16'hffff;
  rom[00325] = 16'hffff;
  rom[00326] = 16'hffff;
  rom[00327] = 16'hffff;
  rom[00328] = 16'hffff;
  rom[00329] = 16'hffff;
  rom[00330] = 16'hffff;
  rom[00331] = 16'hffff;
  rom[00332] = 16'hffff;
  rom[00333] = 16'hffff;
  rom[00334] = 16'hffff;
  rom[00335] = 16'hffff;
  rom[00336] = 16'hffff;
  rom[00337] = 16'hffff;
  rom[00338] = 16'hffff;
  rom[00339] = 16'hffff;
  rom[00340] = 16'hffff;
  rom[00341] = 16'hffff;
  rom[00342] = 16'hffff;
  rom[00343] = 16'hffff;
  rom[00344] = 16'hffff;
  rom[00345] = 16'hffff;
  rom[00346] = 16'hffff;
  rom[00347] = 16'hffff;
  rom[00348] = 16'hffff;
  rom[00349] = 16'hffff;
  rom[00350] = 16'hffff;
  rom[00351] = 16'hffff;
  rom[00352] = 16'hffff;
  rom[00353] = 16'hffff;
  rom[00354] = 16'hffff;
  rom[00355] = 16'hffff;
  rom[00356] = 16'hffff;
  rom[00357] = 16'hffff;
  rom[00358] = 16'hffff;
  rom[00359] = 16'hffff;
  rom[00360] = 16'hffff;
  rom[00361] = 16'hffff;
  rom[00362] = 16'hffff;
  rom[00363] = 16'hffff;
  rom[00364] = 16'hffff;
  rom[00365] = 16'hffff;
  rom[00366] = 16'hffff;
  rom[00367] = 16'hffff;
  rom[00368] = 16'hffff;
  rom[00369] = 16'hffff;
  rom[00370] = 16'hffff;
  rom[00371] = 16'hffff;
  rom[00372] = 16'hffff;
  rom[00373] = 16'hffff;
  rom[00374] = 16'hffff;
  rom[00375] = 16'hffff;
  rom[00376] = 16'hffff;
  rom[00377] = 16'hffff;
  rom[00378] = 16'hffff;
  rom[00379] = 16'hffff;
  rom[00380] = 16'hffff;
  rom[00381] = 16'hffff;
  rom[00382] = 16'hffff;
  rom[00383] = 16'hffff;
  rom[00384] = 16'hffff;
  rom[00385] = 16'hffff;
  rom[00386] = 16'hffff;
  rom[00387] = 16'hffff;
  rom[00388] = 16'hffff;
  rom[00389] = 16'hffff;
  rom[00390] = 16'hffff;
  rom[00391] = 16'hffff;
  rom[00392] = 16'hffff;
  rom[00393] = 16'hffff;
  rom[00394] = 16'hffff;
  rom[00395] = 16'hffff;
  rom[00396] = 16'hffff;
  rom[00397] = 16'hffff;
  rom[00398] = 16'hffff;
  rom[00399] = 16'hffff;
  rom[00400] = 16'hffff;
  rom[00401] = 16'hffff;
  rom[00402] = 16'hffff;
  rom[00403] = 16'hffff;
  rom[00404] = 16'hffff;
  rom[00405] = 16'hffff;
  rom[00406] = 16'hffff;
  rom[00407] = 16'hffff;
  rom[00408] = 16'hffff;
  rom[00409] = 16'hffff;
  rom[00410] = 16'hffff;
  rom[00411] = 16'hffff;
  rom[00412] = 16'hffff;
  rom[00413] = 16'hffff;
  rom[00414] = 16'hffff;
  rom[00415] = 16'hffff;
  rom[00416] = 16'hffff;
  rom[00417] = 16'hffff;
  rom[00418] = 16'hffff;
  rom[00419] = 16'hffff;
  rom[00420] = 16'hffff;
  rom[00421] = 16'hffff;
  rom[00422] = 16'hffff;
  rom[00423] = 16'hffff;
  rom[00424] = 16'hffff;
  rom[00425] = 16'hffff;
  rom[00426] = 16'hffff;
  rom[00427] = 16'hffff;
  rom[00428] = 16'hffff;
  rom[00429] = 16'hffff;
  rom[00430] = 16'hffff;
  rom[00431] = 16'hffff;
  rom[00432] = 16'hffff;
  rom[00433] = 16'hffff;
  rom[00434] = 16'hffff;
  rom[00435] = 16'hffff;
  rom[00436] = 16'hffff;
  rom[00437] = 16'hffff;
  rom[00438] = 16'hffff;
  rom[00439] = 16'hffff;
  rom[00440] = 16'hffff;
  rom[00441] = 16'hffff;
  rom[00442] = 16'hffff;
  rom[00443] = 16'hffff;
  rom[00444] = 16'hffff;
  rom[00445] = 16'hffff;
  rom[00446] = 16'hffff;
  rom[00447] = 16'hffff;
  rom[00448] = 16'hffff;
  rom[00449] = 16'hffff;
  rom[00450] = 16'hffff;
  rom[00451] = 16'hffff;
  rom[00452] = 16'hffff;
  rom[00453] = 16'hffff;
  rom[00454] = 16'hffff;
  rom[00455] = 16'hffff;
  rom[00456] = 16'hffdf;
  rom[00457] = 16'hffff;
  rom[00458] = 16'hffff;
  rom[00459] = 16'hffff;
  rom[00460] = 16'hffff;
  rom[00461] = 16'hffff;
  rom[00462] = 16'hffff;
  rom[00463] = 16'hffff;
  rom[00464] = 16'hffff;
  rom[00465] = 16'hffff;
  rom[00466] = 16'hffff;
  rom[00467] = 16'hffff;
  rom[00468] = 16'hffff;
  rom[00469] = 16'hffff;
  rom[00470] = 16'hffff;
  rom[00471] = 16'hffff;
  rom[00472] = 16'hffff;
  rom[00473] = 16'hffff;
  rom[00474] = 16'hffff;
  rom[00475] = 16'hffff;
  rom[00476] = 16'hffff;
  rom[00477] = 16'hffff;
  rom[00478] = 16'hffff;
  rom[00479] = 16'hffff;
  rom[00480] = 16'hffff;
  rom[00481] = 16'hffff;
  rom[00482] = 16'hffff;
  rom[00483] = 16'hffff;
  rom[00484] = 16'hffff;
  rom[00485] = 16'hffff;
  rom[00486] = 16'hffde;
  rom[00487] = 16'hffff;
  rom[00488] = 16'hfffe;
  rom[00489] = 16'ha4b0;
  rom[00490] = 16'hbc8d;
  rom[00491] = 16'he54e;
  rom[00492] = 16'hdd2d;
  rom[00493] = 16'hdd2d;
  rom[00494] = 16'hd50c;
  rom[00495] = 16'hbc6b;
  rom[00496] = 16'h82e6;
  rom[00497] = 16'h3921;
  rom[00498] = 16'h28c0;
  rom[00499] = 16'h6aea;
  rom[00500] = 16'hf73c;
  rom[00501] = 16'hffff;
  rom[00502] = 16'hffde;
  rom[00503] = 16'hffff;
  rom[00504] = 16'hffff;
  rom[00505] = 16'hffff;
  rom[00506] = 16'hffde;
  rom[00507] = 16'hffff;
  rom[00508] = 16'hffff;
  rom[00509] = 16'hffff;
  rom[00510] = 16'hfffe;
  rom[00511] = 16'hffff;
  rom[00512] = 16'hffdf;
  rom[00513] = 16'hffff;
  rom[00514] = 16'hffff;
  rom[00515] = 16'hffff;
  rom[00516] = 16'hffff;
  rom[00517] = 16'hffff;
  rom[00518] = 16'hffff;
  rom[00519] = 16'hffff;
  rom[00520] = 16'hffff;
  rom[00521] = 16'hffff;
  rom[00522] = 16'hffff;
  rom[00523] = 16'hffff;
  rom[00524] = 16'hffff;
  rom[00525] = 16'hffff;
  rom[00526] = 16'hffff;
  rom[00527] = 16'hffff;
  rom[00528] = 16'hffff;
  rom[00529] = 16'hffff;
  rom[00530] = 16'hffff;
  rom[00531] = 16'hffff;
  rom[00532] = 16'hffff;
  rom[00533] = 16'hffff;
  rom[00534] = 16'hffff;
  rom[00535] = 16'hffff;
  rom[00536] = 16'hffdf;
  rom[00537] = 16'hffff;
  rom[00538] = 16'hffff;
  rom[00539] = 16'hffff;
  rom[00540] = 16'hffff;
  rom[00541] = 16'hffff;
  rom[00542] = 16'hffff;
  rom[00543] = 16'hffff;
  rom[00544] = 16'hffff;
  rom[00545] = 16'hffff;
  rom[00546] = 16'hffff;
  rom[00547] = 16'hffff;
  rom[00548] = 16'hffff;
  rom[00549] = 16'hffff;
  rom[00550] = 16'hffff;
  rom[00551] = 16'hffff;
  rom[00552] = 16'hffff;
  rom[00553] = 16'hffff;
  rom[00554] = 16'hffff;
  rom[00555] = 16'hffff;
  rom[00556] = 16'hffff;
  rom[00557] = 16'hffff;
  rom[00558] = 16'hffff;
  rom[00559] = 16'hffff;
  rom[00560] = 16'hffff;
  rom[00561] = 16'hffff;
  rom[00562] = 16'hffff;
  rom[00563] = 16'hffff;
  rom[00564] = 16'hffff;
  rom[00565] = 16'hffff;
  rom[00566] = 16'hffff;
  rom[00567] = 16'hffff;
  rom[00568] = 16'hffff;
  rom[00569] = 16'hffff;
  rom[00570] = 16'hffff;
  rom[00571] = 16'hffff;
  rom[00572] = 16'hffff;
  rom[00573] = 16'hffff;
  rom[00574] = 16'hffff;
  rom[00575] = 16'hffff;
  rom[00576] = 16'hffff;
  rom[00577] = 16'hffff;
  rom[00578] = 16'hffff;
  rom[00579] = 16'hffff;
  rom[00580] = 16'hffff;
  rom[00581] = 16'hffff;
  rom[00582] = 16'hffff;
  rom[00583] = 16'hffff;
  rom[00584] = 16'hffff;
  rom[00585] = 16'hffff;
  rom[00586] = 16'hffff;
  rom[00587] = 16'hffff;
  rom[00588] = 16'hffff;
  rom[00589] = 16'hffff;
  rom[00590] = 16'hffff;
  rom[00591] = 16'hffff;
  rom[00592] = 16'hffff;
  rom[00593] = 16'hffff;
  rom[00594] = 16'hffff;
  rom[00595] = 16'hffff;
  rom[00596] = 16'hffff;
  rom[00597] = 16'hffff;
  rom[00598] = 16'hffff;
  rom[00599] = 16'hffff;
  rom[00600] = 16'hffff;
  rom[00601] = 16'hffff;
  rom[00602] = 16'hffff;
  rom[00603] = 16'hffff;
  rom[00604] = 16'hffff;
  rom[00605] = 16'hffff;
  rom[00606] = 16'hffff;
  rom[00607] = 16'hffff;
  rom[00608] = 16'hffff;
  rom[00609] = 16'hffff;
  rom[00610] = 16'hffff;
  rom[00611] = 16'hffff;
  rom[00612] = 16'hffff;
  rom[00613] = 16'hffff;
  rom[00614] = 16'hffff;
  rom[00615] = 16'hffff;
  rom[00616] = 16'hffff;
  rom[00617] = 16'hffff;
  rom[00618] = 16'hffff;
  rom[00619] = 16'hffff;
  rom[00620] = 16'hffff;
  rom[00621] = 16'hffff;
  rom[00622] = 16'hffff;
  rom[00623] = 16'hffff;
  rom[00624] = 16'hffff;
  rom[00625] = 16'hffff;
  rom[00626] = 16'hffff;
  rom[00627] = 16'hffff;
  rom[00628] = 16'hffff;
  rom[00629] = 16'hffff;
  rom[00630] = 16'hffff;
  rom[00631] = 16'hffff;
  rom[00632] = 16'hffff;
  rom[00633] = 16'hffff;
  rom[00634] = 16'hffff;
  rom[00635] = 16'hffff;
  rom[00636] = 16'hffff;
  rom[00637] = 16'hffff;
  rom[00638] = 16'hffff;
  rom[00639] = 16'hffff;
  rom[00640] = 16'hffff;
  rom[00641] = 16'hffff;
  rom[00642] = 16'hffff;
  rom[00643] = 16'hffff;
  rom[00644] = 16'hffff;
  rom[00645] = 16'hffff;
  rom[00646] = 16'hffff;
  rom[00647] = 16'hffff;
  rom[00648] = 16'hffff;
  rom[00649] = 16'hffff;
  rom[00650] = 16'hffff;
  rom[00651] = 16'hffff;
  rom[00652] = 16'hffff;
  rom[00653] = 16'hffff;
  rom[00654] = 16'hffff;
  rom[00655] = 16'hffdf;
  rom[00656] = 16'hffff;
  rom[00657] = 16'hffbf;
  rom[00658] = 16'hef5d;
  rom[00659] = 16'hd67a;
  rom[00660] = 16'hce39;
  rom[00661] = 16'hc618;
  rom[00662] = 16'hc5f8;
  rom[00663] = 16'hc638;
  rom[00664] = 16'hdedb;
  rom[00665] = 16'hef3d;
  rom[00666] = 16'hffdf;
  rom[00667] = 16'hffff;
  rom[00668] = 16'hffff;
  rom[00669] = 16'hffff;
  rom[00670] = 16'hffff;
  rom[00671] = 16'hffff;
  rom[00672] = 16'hffff;
  rom[00673] = 16'hffff;
  rom[00674] = 16'hffff;
  rom[00675] = 16'hffff;
  rom[00676] = 16'hffff;
  rom[00677] = 16'hffff;
  rom[00678] = 16'hffff;
  rom[00679] = 16'hffff;
  rom[00680] = 16'hffff;
  rom[00681] = 16'hffff;
  rom[00682] = 16'hffff;
  rom[00683] = 16'hffff;
  rom[00684] = 16'hffff;
  rom[00685] = 16'hffff;
  rom[00686] = 16'hffff;
  rom[00687] = 16'hfffe;
  rom[00688] = 16'hfffe;
  rom[00689] = 16'ha4b0;
  rom[00690] = 16'hcccc;
  rom[00691] = 16'he52a;
  rom[00692] = 16'hfd6c;
  rom[00693] = 16'hed2a;
  rom[00694] = 16'hf54a;
  rom[00695] = 16'hed2a;
  rom[00696] = 16'hdd2c;
  rom[00697] = 16'hbc8b;
  rom[00698] = 16'h82e6;
  rom[00699] = 16'h51a4;
  rom[00700] = 16'hddd7;
  rom[00701] = 16'hff9e;
  rom[00702] = 16'hffff;
  rom[00703] = 16'hffff;
  rom[00704] = 16'hffff;
  rom[00705] = 16'hffff;
  rom[00706] = 16'hffff;
  rom[00707] = 16'hffff;
  rom[00708] = 16'hffff;
  rom[00709] = 16'hffff;
  rom[00710] = 16'hffff;
  rom[00711] = 16'hffff;
  rom[00712] = 16'hffff;
  rom[00713] = 16'hffff;
  rom[00714] = 16'hffff;
  rom[00715] = 16'hffff;
  rom[00716] = 16'hffff;
  rom[00717] = 16'hffff;
  rom[00718] = 16'hffff;
  rom[00719] = 16'hffff;
  rom[00720] = 16'hffff;
  rom[00721] = 16'hffff;
  rom[00722] = 16'hffff;
  rom[00723] = 16'hffff;
  rom[00724] = 16'hffff;
  rom[00725] = 16'hffff;
  rom[00726] = 16'hffdf;
  rom[00727] = 16'hdebb;
  rom[00728] = 16'hb596;
  rom[00729] = 16'h83f0;
  rom[00730] = 16'h630c;
  rom[00731] = 16'h5acb;
  rom[00732] = 16'h526a;
  rom[00733] = 16'h528a;
  rom[00734] = 16'h6b4d;
  rom[00735] = 16'h9492;
  rom[00736] = 16'hc5f8;
  rom[00737] = 16'he71c;
  rom[00738] = 16'hffff;
  rom[00739] = 16'hffff;
  rom[00740] = 16'hffff;
  rom[00741] = 16'hffff;
  rom[00742] = 16'hffff;
  rom[00743] = 16'hffff;
  rom[00744] = 16'hffff;
  rom[00745] = 16'hffff;
  rom[00746] = 16'hffff;
  rom[00747] = 16'hffff;
  rom[00748] = 16'hffff;
  rom[00749] = 16'hffff;
  rom[00750] = 16'hffff;
  rom[00751] = 16'hffff;
  rom[00752] = 16'hffff;
  rom[00753] = 16'hffff;
  rom[00754] = 16'hffff;
  rom[00755] = 16'hffff;
  rom[00756] = 16'hffff;
  rom[00757] = 16'hffff;
  rom[00758] = 16'hffff;
  rom[00759] = 16'hffff;
  rom[00760] = 16'hffff;
  rom[00761] = 16'hffff;
  rom[00762] = 16'hffff;
  rom[00763] = 16'hffff;
  rom[00764] = 16'hffff;
  rom[00765] = 16'hffff;
  rom[00766] = 16'hffff;
  rom[00767] = 16'hffff;
  rom[00768] = 16'hffff;
  rom[00769] = 16'hffff;
  rom[00770] = 16'hffff;
  rom[00771] = 16'hffff;
  rom[00772] = 16'hffff;
  rom[00773] = 16'hffff;
  rom[00774] = 16'hffff;
  rom[00775] = 16'hffff;
  rom[00776] = 16'hffff;
  rom[00777] = 16'hffff;
  rom[00778] = 16'hffff;
  rom[00779] = 16'hffff;
  rom[00780] = 16'hffff;
  rom[00781] = 16'hffff;
  rom[00782] = 16'hffff;
  rom[00783] = 16'hffff;
  rom[00784] = 16'hffff;
  rom[00785] = 16'hffff;
  rom[00786] = 16'hffff;
  rom[00787] = 16'hffff;
  rom[00788] = 16'hffff;
  rom[00789] = 16'hffff;
  rom[00790] = 16'hffff;
  rom[00791] = 16'hffff;
  rom[00792] = 16'hffff;
  rom[00793] = 16'hffff;
  rom[00794] = 16'hffff;
  rom[00795] = 16'hffff;
  rom[00796] = 16'hffff;
  rom[00797] = 16'hffff;
  rom[00798] = 16'hffff;
  rom[00799] = 16'hffff;
  rom[00800] = 16'hffff;
  rom[00801] = 16'hffff;
  rom[00802] = 16'hffff;
  rom[00803] = 16'hffff;
  rom[00804] = 16'hffff;
  rom[00805] = 16'hffff;
  rom[00806] = 16'hffff;
  rom[00807] = 16'hffff;
  rom[00808] = 16'hffff;
  rom[00809] = 16'hffff;
  rom[00810] = 16'hffff;
  rom[00811] = 16'hffff;
  rom[00812] = 16'hffff;
  rom[00813] = 16'hffff;
  rom[00814] = 16'hffff;
  rom[00815] = 16'hffff;
  rom[00816] = 16'hffff;
  rom[00817] = 16'hffff;
  rom[00818] = 16'hffff;
  rom[00819] = 16'hffff;
  rom[00820] = 16'hffff;
  rom[00821] = 16'hffff;
  rom[00822] = 16'hffff;
  rom[00823] = 16'hffff;
  rom[00824] = 16'hffff;
  rom[00825] = 16'hffff;
  rom[00826] = 16'hffff;
  rom[00827] = 16'hffff;
  rom[00828] = 16'hffff;
  rom[00829] = 16'hffff;
  rom[00830] = 16'hffff;
  rom[00831] = 16'hffff;
  rom[00832] = 16'hffff;
  rom[00833] = 16'hffff;
  rom[00834] = 16'hffff;
  rom[00835] = 16'hffff;
  rom[00836] = 16'hffff;
  rom[00837] = 16'hffff;
  rom[00838] = 16'hffff;
  rom[00839] = 16'hffff;
  rom[00840] = 16'hffff;
  rom[00841] = 16'hffff;
  rom[00842] = 16'hffff;
  rom[00843] = 16'hffff;
  rom[00844] = 16'hffff;
  rom[00845] = 16'hffff;
  rom[00846] = 16'hffff;
  rom[00847] = 16'hffff;
  rom[00848] = 16'hffff;
  rom[00849] = 16'hffff;
  rom[00850] = 16'hffff;
  rom[00851] = 16'hffff;
  rom[00852] = 16'hffff;
  rom[00853] = 16'hffff;
  rom[00854] = 16'hffff;
  rom[00855] = 16'hffbe;
  rom[00856] = 16'hce59;
  rom[00857] = 16'h7baf;
  rom[00858] = 16'h4228;
  rom[00859] = 16'h3186;
  rom[00860] = 16'h18e3;
  rom[00861] = 16'h18c3;
  rom[00862] = 16'h1082;
  rom[00863] = 16'h20e4;
  rom[00864] = 16'h39c7;
  rom[00865] = 16'h4a49;
  rom[00866] = 16'h7bcf;
  rom[00867] = 16'hd6ba;
  rom[00868] = 16'hffdf;
  rom[00869] = 16'hffff;
  rom[00870] = 16'hffff;
  rom[00871] = 16'hffff;
  rom[00872] = 16'hffff;
  rom[00873] = 16'hffff;
  rom[00874] = 16'hffff;
  rom[00875] = 16'hffff;
  rom[00876] = 16'hffff;
  rom[00877] = 16'hffff;
  rom[00878] = 16'hffff;
  rom[00879] = 16'hffff;
  rom[00880] = 16'hffff;
  rom[00881] = 16'hffff;
  rom[00882] = 16'hffff;
  rom[00883] = 16'hffff;
  rom[00884] = 16'hffff;
  rom[00885] = 16'hffff;
  rom[00886] = 16'hffff;
  rom[00887] = 16'hffff;
  rom[00888] = 16'hffde;
  rom[00889] = 16'h9caf;
  rom[00890] = 16'hc489;
  rom[00891] = 16'hfd49;
  rom[00892] = 16'hfd48;
  rom[00893] = 16'hfd49;
  rom[00894] = 16'hf507;
  rom[00895] = 16'hfd49;
  rom[00896] = 16'hed29;
  rom[00897] = 16'hed6c;
  rom[00898] = 16'hd4ec;
  rom[00899] = 16'habea;
  rom[00900] = 16'h7226;
  rom[00901] = 16'hcd53;
  rom[00902] = 16'hff9d;
  rom[00903] = 16'hffff;
  rom[00904] = 16'hffff;
  rom[00905] = 16'hffff;
  rom[00906] = 16'hffff;
  rom[00907] = 16'hffff;
  rom[00908] = 16'hffff;
  rom[00909] = 16'hffff;
  rom[00910] = 16'hffff;
  rom[00911] = 16'hffff;
  rom[00912] = 16'hffdf;
  rom[00913] = 16'hffff;
  rom[00914] = 16'hffff;
  rom[00915] = 16'hffff;
  rom[00916] = 16'hffff;
  rom[00917] = 16'hffff;
  rom[00918] = 16'hffff;
  rom[00919] = 16'hffff;
  rom[00920] = 16'hffff;
  rom[00921] = 16'hffff;
  rom[00922] = 16'hffff;
  rom[00923] = 16'hffff;
  rom[00924] = 16'hffdf;
  rom[00925] = 16'hef1c;
  rom[00926] = 16'h8c30;
  rom[00927] = 16'h3145;
  rom[00928] = 16'h18e3;
  rom[00929] = 16'h18c3;
  rom[00930] = 16'h1082;
  rom[00931] = 16'h18a3;
  rom[00932] = 16'h10c2;
  rom[00933] = 16'h18e3;
  rom[00934] = 16'h1082;
  rom[00935] = 16'h18c3;
  rom[00936] = 16'h1903;
  rom[00937] = 16'h4a69;
  rom[00938] = 16'ha534;
  rom[00939] = 16'hf77e;
  rom[00940] = 16'hffff;
  rom[00941] = 16'hffff;
  rom[00942] = 16'hffff;
  rom[00943] = 16'hffff;
  rom[00944] = 16'hffff;
  rom[00945] = 16'hffff;
  rom[00946] = 16'hffff;
  rom[00947] = 16'hffff;
  rom[00948] = 16'hffff;
  rom[00949] = 16'hffff;
  rom[00950] = 16'hffff;
  rom[00951] = 16'hffff;
  rom[00952] = 16'hffff;
  rom[00953] = 16'hffff;
  rom[00954] = 16'hffff;
  rom[00955] = 16'hffff;
  rom[00956] = 16'hffff;
  rom[00957] = 16'hffff;
  rom[00958] = 16'hffff;
  rom[00959] = 16'hffff;
  rom[00960] = 16'hffff;
  rom[00961] = 16'hffff;
  rom[00962] = 16'hffff;
  rom[00963] = 16'hffff;
  rom[00964] = 16'hffff;
  rom[00965] = 16'hffff;
  rom[00966] = 16'hffff;
  rom[00967] = 16'hffff;
  rom[00968] = 16'hffff;
  rom[00969] = 16'hffff;
  rom[00970] = 16'hffff;
  rom[00971] = 16'hffff;
  rom[00972] = 16'hffff;
  rom[00973] = 16'hffff;
  rom[00974] = 16'hffff;
  rom[00975] = 16'hffff;
  rom[00976] = 16'hffff;
  rom[00977] = 16'hffff;
  rom[00978] = 16'hffff;
  rom[00979] = 16'hffff;
  rom[00980] = 16'hffff;
  rom[00981] = 16'hffff;
  rom[00982] = 16'hffff;
  rom[00983] = 16'hffff;
  rom[00984] = 16'hffff;
  rom[00985] = 16'hffff;
  rom[00986] = 16'hffff;
  rom[00987] = 16'hffff;
  rom[00988] = 16'hffff;
  rom[00989] = 16'hffff;
  rom[00990] = 16'hffff;
  rom[00991] = 16'hffff;
  rom[00992] = 16'hffff;
  rom[00993] = 16'hffff;
  rom[00994] = 16'hffff;
  rom[00995] = 16'hffff;
  rom[00996] = 16'hffff;
  rom[00997] = 16'hffff;
  rom[00998] = 16'hffff;
  rom[00999] = 16'hffff;
  rom[01000] = 16'hffff;
  rom[01001] = 16'hffff;
  rom[01002] = 16'hffff;
  rom[01003] = 16'hffff;
  rom[01004] = 16'hffff;
  rom[01005] = 16'hffff;
  rom[01006] = 16'hffff;
  rom[01007] = 16'hffff;
  rom[01008] = 16'hffff;
  rom[01009] = 16'hffff;
  rom[01010] = 16'hffff;
  rom[01011] = 16'hffff;
  rom[01012] = 16'hffff;
  rom[01013] = 16'hffff;
  rom[01014] = 16'hffff;
  rom[01015] = 16'hffff;
  rom[01016] = 16'hffff;
  rom[01017] = 16'hffff;
  rom[01018] = 16'hffff;
  rom[01019] = 16'hffff;
  rom[01020] = 16'hffff;
  rom[01021] = 16'hffff;
  rom[01022] = 16'hffff;
  rom[01023] = 16'hffff;
  rom[01024] = 16'hffff;
  rom[01025] = 16'hffff;
  rom[01026] = 16'hffff;
  rom[01027] = 16'hffff;
  rom[01028] = 16'hffff;
  rom[01029] = 16'hffff;
  rom[01030] = 16'hffff;
  rom[01031] = 16'hffff;
  rom[01032] = 16'hffff;
  rom[01033] = 16'hffff;
  rom[01034] = 16'hffff;
  rom[01035] = 16'hffff;
  rom[01036] = 16'hffff;
  rom[01037] = 16'hffff;
  rom[01038] = 16'hffff;
  rom[01039] = 16'hffff;
  rom[01040] = 16'hffff;
  rom[01041] = 16'hffff;
  rom[01042] = 16'hffff;
  rom[01043] = 16'hffff;
  rom[01044] = 16'hffff;
  rom[01045] = 16'hffff;
  rom[01046] = 16'hffff;
  rom[01047] = 16'hffff;
  rom[01048] = 16'hffff;
  rom[01049] = 16'hffff;
  rom[01050] = 16'hffff;
  rom[01051] = 16'hffff;
  rom[01052] = 16'hffff;
  rom[01053] = 16'hffff;
  rom[01054] = 16'hffdf;
  rom[01055] = 16'h9cd3;
  rom[01056] = 16'h3186;
  rom[01057] = 16'h0861;
  rom[01058] = 16'h18c3;
  rom[01059] = 16'h1082;
  rom[01060] = 16'h10a2;
  rom[01061] = 16'h10a2;
  rom[01062] = 16'h2104;
  rom[01063] = 16'h18c3;
  rom[01064] = 16'h1082;
  rom[01065] = 16'h10c2;
  rom[01066] = 16'h18c3;
  rom[01067] = 16'h2965;
  rom[01068] = 16'had75;
  rom[01069] = 16'hffdf;
  rom[01070] = 16'hffff;
  rom[01071] = 16'hffdf;
  rom[01072] = 16'hffff;
  rom[01073] = 16'hffff;
  rom[01074] = 16'hffff;
  rom[01075] = 16'hffff;
  rom[01076] = 16'hffff;
  rom[01077] = 16'hffff;
  rom[01078] = 16'hffff;
  rom[01079] = 16'hffff;
  rom[01080] = 16'hffff;
  rom[01081] = 16'hffff;
  rom[01082] = 16'hffff;
  rom[01083] = 16'hffff;
  rom[01084] = 16'hffff;
  rom[01085] = 16'hffff;
  rom[01086] = 16'hffff;
  rom[01087] = 16'hffff;
  rom[01088] = 16'hffff;
  rom[01089] = 16'h9caf;
  rom[01090] = 16'hccca;
  rom[01091] = 16'hf527;
  rom[01092] = 16'hfd27;
  rom[01093] = 16'hfd27;
  rom[01094] = 16'hfd47;
  rom[01095] = 16'hfd27;
  rom[01096] = 16'hfd69;
  rom[01097] = 16'he4e8;
  rom[01098] = 16'hfdad;
  rom[01099] = 16'hdd0c;
  rom[01100] = 16'hd4ed;
  rom[01101] = 16'h7aa5;
  rom[01102] = 16'hbd11;
  rom[01103] = 16'hffbd;
  rom[01104] = 16'hf7df;
  rom[01105] = 16'hf7df;
  rom[01106] = 16'hffff;
  rom[01107] = 16'hffbf;
  rom[01108] = 16'hffff;
  rom[01109] = 16'hffff;
  rom[01110] = 16'hffff;
  rom[01111] = 16'hffff;
  rom[01112] = 16'hffff;
  rom[01113] = 16'hffff;
  rom[01114] = 16'hffff;
  rom[01115] = 16'hffff;
  rom[01116] = 16'hffff;
  rom[01117] = 16'hffff;
  rom[01118] = 16'hffff;
  rom[01119] = 16'hffff;
  rom[01120] = 16'hffff;
  rom[01121] = 16'hffff;
  rom[01122] = 16'hffff;
  rom[01123] = 16'hffff;
  rom[01124] = 16'hef1c;
  rom[01125] = 16'h528a;
  rom[01126] = 16'h18a3;
  rom[01127] = 16'h1882;
  rom[01128] = 16'h18c3;
  rom[01129] = 16'h0861;
  rom[01130] = 16'h18e3;
  rom[01131] = 16'h18c3;
  rom[01132] = 16'h18c3;
  rom[01133] = 16'h0861;
  rom[01134] = 16'h18a3;
  rom[01135] = 16'h10a2;
  rom[01136] = 16'h10a2;
  rom[01137] = 16'h10a2;
  rom[01138] = 16'h2104;
  rom[01139] = 16'h9471;
  rom[01140] = 16'hffbf;
  rom[01141] = 16'hffff;
  rom[01142] = 16'hffff;
  rom[01143] = 16'hffff;
  rom[01144] = 16'hffff;
  rom[01145] = 16'hffff;
  rom[01146] = 16'hffff;
  rom[01147] = 16'hffff;
  rom[01148] = 16'hffff;
  rom[01149] = 16'hffff;
  rom[01150] = 16'hffff;
  rom[01151] = 16'hffff;
  rom[01152] = 16'hffff;
  rom[01153] = 16'hffff;
  rom[01154] = 16'hffff;
  rom[01155] = 16'hffff;
  rom[01156] = 16'hffff;
  rom[01157] = 16'hffff;
  rom[01158] = 16'hffff;
  rom[01159] = 16'hffff;
  rom[01160] = 16'hffff;
  rom[01161] = 16'hffff;
  rom[01162] = 16'hffff;
  rom[01163] = 16'hffff;
  rom[01164] = 16'hffff;
  rom[01165] = 16'hffff;
  rom[01166] = 16'hffff;
  rom[01167] = 16'hffff;
  rom[01168] = 16'hffff;
  rom[01169] = 16'hffff;
  rom[01170] = 16'hffff;
  rom[01171] = 16'hffff;
  rom[01172] = 16'hffff;
  rom[01173] = 16'hffff;
  rom[01174] = 16'hffff;
  rom[01175] = 16'hffff;
  rom[01176] = 16'hffff;
  rom[01177] = 16'hffff;
  rom[01178] = 16'hffff;
  rom[01179] = 16'hffff;
  rom[01180] = 16'hffff;
  rom[01181] = 16'hffff;
  rom[01182] = 16'hffff;
  rom[01183] = 16'hffff;
  rom[01184] = 16'hffff;
  rom[01185] = 16'hffff;
  rom[01186] = 16'hffff;
  rom[01187] = 16'hffff;
  rom[01188] = 16'hffff;
  rom[01189] = 16'hffff;
  rom[01190] = 16'hffff;
  rom[01191] = 16'hffff;
  rom[01192] = 16'hffff;
  rom[01193] = 16'hffff;
  rom[01194] = 16'hffff;
  rom[01195] = 16'hffff;
  rom[01196] = 16'hffff;
  rom[01197] = 16'hffff;
  rom[01198] = 16'hffff;
  rom[01199] = 16'hffff;
  rom[01200] = 16'hffff;
  rom[01201] = 16'hffff;
  rom[01202] = 16'hffff;
  rom[01203] = 16'hffff;
  rom[01204] = 16'hffff;
  rom[01205] = 16'hffff;
  rom[01206] = 16'hffff;
  rom[01207] = 16'hffff;
  rom[01208] = 16'hffff;
  rom[01209] = 16'hffff;
  rom[01210] = 16'hffff;
  rom[01211] = 16'hffff;
  rom[01212] = 16'hffff;
  rom[01213] = 16'hffff;
  rom[01214] = 16'hffff;
  rom[01215] = 16'hffff;
  rom[01216] = 16'hffff;
  rom[01217] = 16'hffff;
  rom[01218] = 16'hffff;
  rom[01219] = 16'hffff;
  rom[01220] = 16'hffff;
  rom[01221] = 16'hffff;
  rom[01222] = 16'hffff;
  rom[01223] = 16'hffff;
  rom[01224] = 16'hffff;
  rom[01225] = 16'hffff;
  rom[01226] = 16'hffff;
  rom[01227] = 16'hffff;
  rom[01228] = 16'hffff;
  rom[01229] = 16'hffff;
  rom[01230] = 16'hffff;
  rom[01231] = 16'hffff;
  rom[01232] = 16'hffff;
  rom[01233] = 16'hffff;
  rom[01234] = 16'hffff;
  rom[01235] = 16'hffff;
  rom[01236] = 16'hffff;
  rom[01237] = 16'hffff;
  rom[01238] = 16'hffff;
  rom[01239] = 16'hffff;
  rom[01240] = 16'hffff;
  rom[01241] = 16'hffff;
  rom[01242] = 16'hffff;
  rom[01243] = 16'hffff;
  rom[01244] = 16'hffff;
  rom[01245] = 16'hffff;
  rom[01246] = 16'hffff;
  rom[01247] = 16'hffff;
  rom[01248] = 16'hffff;
  rom[01249] = 16'hffff;
  rom[01250] = 16'hffff;
  rom[01251] = 16'hffff;
  rom[01252] = 16'hffdf;
  rom[01253] = 16'hffbf;
  rom[01254] = 16'h9492;
  rom[01255] = 16'h2144;
  rom[01256] = 16'h1081;
  rom[01257] = 16'h18c3;
  rom[01258] = 16'h10a2;
  rom[01259] = 16'h18e3;
  rom[01260] = 16'h10c2;
  rom[01261] = 16'h18a3;
  rom[01262] = 16'h1082;
  rom[01263] = 16'h10a2;
  rom[01264] = 16'h18c3;
  rom[01265] = 16'h18e3;
  rom[01266] = 16'h10a2;
  rom[01267] = 16'h10a2;
  rom[01268] = 16'h31a6;
  rom[01269] = 16'hbdb6;
  rom[01270] = 16'hf7be;
  rom[01271] = 16'hffff;
  rom[01272] = 16'hffff;
  rom[01273] = 16'hffff;
  rom[01274] = 16'hffff;
  rom[01275] = 16'hffff;
  rom[01276] = 16'hffff;
  rom[01277] = 16'hffff;
  rom[01278] = 16'hffff;
  rom[01279] = 16'hffff;
  rom[01280] = 16'hffbf;
  rom[01281] = 16'hef5d;
  rom[01282] = 16'hf79d;
  rom[01283] = 16'hfffe;
  rom[01284] = 16'hfffe;
  rom[01285] = 16'hffff;
  rom[01286] = 16'hffff;
  rom[01287] = 16'hffff;
  rom[01288] = 16'hffff;
  rom[01289] = 16'h9cb0;
  rom[01290] = 16'hc489;
  rom[01291] = 16'hfd68;
  rom[01292] = 16'hfd28;
  rom[01293] = 16'hfd28;
  rom[01294] = 16'hfd27;
  rom[01295] = 16'hfd28;
  rom[01296] = 16'hfd28;
  rom[01297] = 16'hfd6a;
  rom[01298] = 16'he508;
  rom[01299] = 16'hf56b;
  rom[01300] = 16'hed2a;
  rom[01301] = 16'hcc8a;
  rom[01302] = 16'h7284;
  rom[01303] = 16'ha46d;
  rom[01304] = 16'hf79c;
  rom[01305] = 16'hffff;
  rom[01306] = 16'hffdf;
  rom[01307] = 16'hffff;
  rom[01308] = 16'hd679;
  rom[01309] = 16'hb554;
  rom[01310] = 16'hd677;
  rom[01311] = 16'hffbd;
  rom[01312] = 16'hffdf;
  rom[01313] = 16'hffff;
  rom[01314] = 16'hffdf;
  rom[01315] = 16'hffff;
  rom[01316] = 16'hffff;
  rom[01317] = 16'hffff;
  rom[01318] = 16'hffff;
  rom[01319] = 16'hffff;
  rom[01320] = 16'hffdf;
  rom[01321] = 16'hffff;
  rom[01322] = 16'hffff;
  rom[01323] = 16'hef5d;
  rom[01324] = 16'h83ae;
  rom[01325] = 16'h18a3;
  rom[01326] = 16'h10a2;
  rom[01327] = 16'h18c2;
  rom[01328] = 16'h1082;
  rom[01329] = 16'h18c3;
  rom[01330] = 16'h10a2;
  rom[01331] = 16'h10a2;
  rom[01332] = 16'h1082;
  rom[01333] = 16'h18c3;
  rom[01334] = 16'h10a2;
  rom[01335] = 16'h18c3;
  rom[01336] = 16'h1081;
  rom[01337] = 16'h10a2;
  rom[01338] = 16'h0861;
  rom[01339] = 16'h31a6;
  rom[01340] = 16'had34;
  rom[01341] = 16'hffff;
  rom[01342] = 16'hffff;
  rom[01343] = 16'hffff;
  rom[01344] = 16'hffff;
  rom[01345] = 16'hffff;
  rom[01346] = 16'hffff;
  rom[01347] = 16'hffff;
  rom[01348] = 16'hffff;
  rom[01349] = 16'hffff;
  rom[01350] = 16'hffff;
  rom[01351] = 16'hffff;
  rom[01352] = 16'hffff;
  rom[01353] = 16'hffff;
  rom[01354] = 16'hffff;
  rom[01355] = 16'hffff;
  rom[01356] = 16'hffff;
  rom[01357] = 16'hffff;
  rom[01358] = 16'hffff;
  rom[01359] = 16'hffff;
  rom[01360] = 16'hffff;
  rom[01361] = 16'hffff;
  rom[01362] = 16'hffff;
  rom[01363] = 16'hffff;
  rom[01364] = 16'hffff;
  rom[01365] = 16'hffff;
  rom[01366] = 16'hffff;
  rom[01367] = 16'hffff;
  rom[01368] = 16'hffff;
  rom[01369] = 16'hffff;
  rom[01370] = 16'hffff;
  rom[01371] = 16'hffff;
  rom[01372] = 16'hffff;
  rom[01373] = 16'hffff;
  rom[01374] = 16'hffff;
  rom[01375] = 16'hffff;
  rom[01376] = 16'hffff;
  rom[01377] = 16'hffff;
  rom[01378] = 16'hffff;
  rom[01379] = 16'hffff;
  rom[01380] = 16'hffff;
  rom[01381] = 16'hffff;
  rom[01382] = 16'hffff;
  rom[01383] = 16'hffff;
  rom[01384] = 16'hffff;
  rom[01385] = 16'hffff;
  rom[01386] = 16'hffff;
  rom[01387] = 16'hffff;
  rom[01388] = 16'hffff;
  rom[01389] = 16'hffff;
  rom[01390] = 16'hffff;
  rom[01391] = 16'hffff;
  rom[01392] = 16'hffff;
  rom[01393] = 16'hffff;
  rom[01394] = 16'hffff;
  rom[01395] = 16'hffff;
  rom[01396] = 16'hffff;
  rom[01397] = 16'hffff;
  rom[01398] = 16'hffff;
  rom[01399] = 16'hffff;
  rom[01400] = 16'hffff;
  rom[01401] = 16'hffff;
  rom[01402] = 16'hffff;
  rom[01403] = 16'hffff;
  rom[01404] = 16'hffff;
  rom[01405] = 16'hffff;
  rom[01406] = 16'hffff;
  rom[01407] = 16'hffff;
  rom[01408] = 16'hffff;
  rom[01409] = 16'hffff;
  rom[01410] = 16'hffff;
  rom[01411] = 16'hffff;
  rom[01412] = 16'hffff;
  rom[01413] = 16'hffff;
  rom[01414] = 16'hffff;
  rom[01415] = 16'hffff;
  rom[01416] = 16'hffff;
  rom[01417] = 16'hffff;
  rom[01418] = 16'hffff;
  rom[01419] = 16'hffff;
  rom[01420] = 16'hffff;
  rom[01421] = 16'hffff;
  rom[01422] = 16'hffff;
  rom[01423] = 16'hffff;
  rom[01424] = 16'hffff;
  rom[01425] = 16'hffff;
  rom[01426] = 16'hffff;
  rom[01427] = 16'hffff;
  rom[01428] = 16'hffff;
  rom[01429] = 16'hffff;
  rom[01430] = 16'hffff;
  rom[01431] = 16'hffff;
  rom[01432] = 16'hffff;
  rom[01433] = 16'hffff;
  rom[01434] = 16'hffff;
  rom[01435] = 16'hffff;
  rom[01436] = 16'hffff;
  rom[01437] = 16'hffff;
  rom[01438] = 16'hffff;
  rom[01439] = 16'hffff;
  rom[01440] = 16'hffff;
  rom[01441] = 16'hffff;
  rom[01442] = 16'hffff;
  rom[01443] = 16'hffff;
  rom[01444] = 16'hffff;
  rom[01445] = 16'hffff;
  rom[01446] = 16'hffff;
  rom[01447] = 16'hffff;
  rom[01448] = 16'hffff;
  rom[01449] = 16'hffff;
  rom[01450] = 16'hffff;
  rom[01451] = 16'hffff;
  rom[01452] = 16'hffff;
  rom[01453] = 16'hce58;
  rom[01454] = 16'h39e7;
  rom[01455] = 16'h10a2;
  rom[01456] = 16'h18e3;
  rom[01457] = 16'h18e3;
  rom[01458] = 16'h18c3;
  rom[01459] = 16'h18c3;
  rom[01460] = 16'h18e3;
  rom[01461] = 16'h18e3;
  rom[01462] = 16'h10c2;
  rom[01463] = 16'h2104;
  rom[01464] = 16'h1062;
  rom[01465] = 16'h0861;
  rom[01466] = 16'h2104;
  rom[01467] = 16'h10a2;
  rom[01468] = 16'h2104;
  rom[01469] = 16'h41e8;
  rom[01470] = 16'hdedb;
  rom[01471] = 16'hffff;
  rom[01472] = 16'hffff;
  rom[01473] = 16'hffff;
  rom[01474] = 16'hffff;
  rom[01475] = 16'hffff;
  rom[01476] = 16'hffff;
  rom[01477] = 16'hffff;
  rom[01478] = 16'hffff;
  rom[01479] = 16'hffdf;
  rom[01480] = 16'hb576;
  rom[01481] = 16'h736d;
  rom[01482] = 16'h9cb1;
  rom[01483] = 16'hef19;
  rom[01484] = 16'hfffd;
  rom[01485] = 16'hffff;
  rom[01486] = 16'hffff;
  rom[01487] = 16'hffff;
  rom[01488] = 16'hffff;
  rom[01489] = 16'h9cb0;
  rom[01490] = 16'hccea;
  rom[01491] = 16'hf548;
  rom[01492] = 16'hfd69;
  rom[01493] = 16'hfd49;
  rom[01494] = 16'hfd49;
  rom[01495] = 16'hfd08;
  rom[01496] = 16'hfd6a;
  rom[01497] = 16'hf548;
  rom[01498] = 16'hfd6a;
  rom[01499] = 16'hf528;
  rom[01500] = 16'hf549;
  rom[01501] = 16'hed4a;
  rom[01502] = 16'hdd4d;
  rom[01503] = 16'h6a43;
  rom[01504] = 16'hb511;
  rom[01505] = 16'hfffe;
  rom[01506] = 16'hffff;
  rom[01507] = 16'hffdf;
  rom[01508] = 16'hc575;
  rom[01509] = 16'h6267;
  rom[01510] = 16'h5a65;
  rom[01511] = 16'had11;
  rom[01512] = 16'hff9e;
  rom[01513] = 16'hffff;
  rom[01514] = 16'hffff;
  rom[01515] = 16'hffdf;
  rom[01516] = 16'hffff;
  rom[01517] = 16'hffff;
  rom[01518] = 16'hffff;
  rom[01519] = 16'hffff;
  rom[01520] = 16'hffdf;
  rom[01521] = 16'hffff;
  rom[01522] = 16'hffff;
  rom[01523] = 16'hbdf7;
  rom[01524] = 16'h2925;
  rom[01525] = 16'h20c3;
  rom[01526] = 16'h10a2;
  rom[01527] = 16'h18c2;
  rom[01528] = 16'h2925;
  rom[01529] = 16'h0841;
  rom[01530] = 16'h10a2;
  rom[01531] = 16'h18c3;
  rom[01532] = 16'h10a2;
  rom[01533] = 16'h10a2;
  rom[01534] = 16'h18e3;
  rom[01535] = 16'h18c2;
  rom[01536] = 16'h1082;
  rom[01537] = 16'h2104;
  rom[01538] = 16'h10a2;
  rom[01539] = 16'h10a2;
  rom[01540] = 16'h62ec;
  rom[01541] = 16'he71c;
  rom[01542] = 16'hffff;
  rom[01543] = 16'hffff;
  rom[01544] = 16'hffff;
  rom[01545] = 16'hffff;
  rom[01546] = 16'hffff;
  rom[01547] = 16'hffff;
  rom[01548] = 16'hffff;
  rom[01549] = 16'hffff;
  rom[01550] = 16'hffff;
  rom[01551] = 16'hffff;
  rom[01552] = 16'hffff;
  rom[01553] = 16'hffff;
  rom[01554] = 16'hffff;
  rom[01555] = 16'hffff;
  rom[01556] = 16'hffff;
  rom[01557] = 16'hffff;
  rom[01558] = 16'hffff;
  rom[01559] = 16'hffff;
  rom[01560] = 16'hffff;
  rom[01561] = 16'hffff;
  rom[01562] = 16'hffff;
  rom[01563] = 16'hffff;
  rom[01564] = 16'hffff;
  rom[01565] = 16'hffff;
  rom[01566] = 16'hffff;
  rom[01567] = 16'hffff;
  rom[01568] = 16'hffff;
  rom[01569] = 16'hffff;
  rom[01570] = 16'hffff;
  rom[01571] = 16'hffff;
  rom[01572] = 16'hffff;
  rom[01573] = 16'hffff;
  rom[01574] = 16'hffff;
  rom[01575] = 16'hffff;
  rom[01576] = 16'hffff;
  rom[01577] = 16'hffff;
  rom[01578] = 16'hffff;
  rom[01579] = 16'hffff;
  rom[01580] = 16'hffff;
  rom[01581] = 16'hffff;
  rom[01582] = 16'hffff;
  rom[01583] = 16'hffff;
  rom[01584] = 16'hffff;
  rom[01585] = 16'hffff;
  rom[01586] = 16'hffff;
  rom[01587] = 16'hffff;
  rom[01588] = 16'hffff;
  rom[01589] = 16'hffff;
  rom[01590] = 16'hffff;
  rom[01591] = 16'hffff;
  rom[01592] = 16'hffff;
  rom[01593] = 16'hffff;
  rom[01594] = 16'hffff;
  rom[01595] = 16'hffff;
  rom[01596] = 16'hffff;
  rom[01597] = 16'hffff;
  rom[01598] = 16'hffff;
  rom[01599] = 16'hffff;
  rom[01600] = 16'hffff;
  rom[01601] = 16'hffff;
  rom[01602] = 16'hffff;
  rom[01603] = 16'hffff;
  rom[01604] = 16'hffff;
  rom[01605] = 16'hffff;
  rom[01606] = 16'hffff;
  rom[01607] = 16'hffff;
  rom[01608] = 16'hffff;
  rom[01609] = 16'hffff;
  rom[01610] = 16'hffff;
  rom[01611] = 16'hffff;
  rom[01612] = 16'hffff;
  rom[01613] = 16'hffff;
  rom[01614] = 16'hffff;
  rom[01615] = 16'hffff;
  rom[01616] = 16'hffff;
  rom[01617] = 16'hffff;
  rom[01618] = 16'hffff;
  rom[01619] = 16'hffff;
  rom[01620] = 16'hffff;
  rom[01621] = 16'hffff;
  rom[01622] = 16'hffff;
  rom[01623] = 16'hffff;
  rom[01624] = 16'hffff;
  rom[01625] = 16'hffff;
  rom[01626] = 16'hffff;
  rom[01627] = 16'hffff;
  rom[01628] = 16'hffff;
  rom[01629] = 16'hffff;
  rom[01630] = 16'hffff;
  rom[01631] = 16'hffff;
  rom[01632] = 16'hffff;
  rom[01633] = 16'hffff;
  rom[01634] = 16'hffff;
  rom[01635] = 16'hffff;
  rom[01636] = 16'hffff;
  rom[01637] = 16'hffff;
  rom[01638] = 16'hffff;
  rom[01639] = 16'hffff;
  rom[01640] = 16'hffff;
  rom[01641] = 16'hffff;
  rom[01642] = 16'hffff;
  rom[01643] = 16'hffff;
  rom[01644] = 16'hffff;
  rom[01645] = 16'hffff;
  rom[01646] = 16'hffff;
  rom[01647] = 16'hffff;
  rom[01648] = 16'hffff;
  rom[01649] = 16'hffff;
  rom[01650] = 16'hffff;
  rom[01651] = 16'hffff;
  rom[01652] = 16'hffdf;
  rom[01653] = 16'h8430;
  rom[01654] = 16'h10a2;
  rom[01655] = 16'h10a2;
  rom[01656] = 16'h10a2;
  rom[01657] = 16'h10a2;
  rom[01658] = 16'h10a2;
  rom[01659] = 16'h18a3;
  rom[01660] = 16'h10a2;
  rom[01661] = 16'h10a2;
  rom[01662] = 16'h10a2;
  rom[01663] = 16'h18a3;
  rom[01664] = 16'h10c2;
  rom[01665] = 16'h18c3;
  rom[01666] = 16'h1082;
  rom[01667] = 16'h18c3;
  rom[01668] = 16'h10a1;
  rom[01669] = 16'h18e3;
  rom[01670] = 16'ha534;
  rom[01671] = 16'hffff;
  rom[01672] = 16'hffff;
  rom[01673] = 16'hffff;
  rom[01674] = 16'hffff;
  rom[01675] = 16'hffff;
  rom[01676] = 16'hffff;
  rom[01677] = 16'hffff;
  rom[01678] = 16'hffff;
  rom[01679] = 16'hffff;
  rom[01680] = 16'hc618;
  rom[01681] = 16'h41c6;
  rom[01682] = 16'h6aea;
  rom[01683] = 16'h83ab;
  rom[01684] = 16'hcdf3;
  rom[01685] = 16'hffbc;
  rom[01686] = 16'hffdf;
  rom[01687] = 16'hffff;
  rom[01688] = 16'hffff;
  rom[01689] = 16'h9c90;
  rom[01690] = 16'hc4ca;
  rom[01691] = 16'hf549;
  rom[01692] = 16'hed49;
  rom[01693] = 16'hfd69;
  rom[01694] = 16'hfd28;
  rom[01695] = 16'hfd48;
  rom[01696] = 16'hf527;
  rom[01697] = 16'hf548;
  rom[01698] = 16'hf548;
  rom[01699] = 16'hfd48;
  rom[01700] = 16'hfd68;
  rom[01701] = 16'hf549;
  rom[01702] = 16'he52a;
  rom[01703] = 16'hcccb;
  rom[01704] = 16'h72c5;
  rom[01705] = 16'hcdf4;
  rom[01706] = 16'hffbd;
  rom[01707] = 16'hffde;
  rom[01708] = 16'hac6f;
  rom[01709] = 16'hb44c;
  rom[01710] = 16'hc4ed;
  rom[01711] = 16'h8b68;
  rom[01712] = 16'h9c8f;
  rom[01713] = 16'hf79d;
  rom[01714] = 16'hffff;
  rom[01715] = 16'hffff;
  rom[01716] = 16'hffdf;
  rom[01717] = 16'hffff;
  rom[01718] = 16'hffff;
  rom[01719] = 16'hffbe;
  rom[01720] = 16'hffff;
  rom[01721] = 16'hffff;
  rom[01722] = 16'hf79e;
  rom[01723] = 16'h9cb3;
  rom[01724] = 16'h18c3;
  rom[01725] = 16'h1082;
  rom[01726] = 16'h10c2;
  rom[01727] = 16'h18a3;
  rom[01728] = 16'h10a2;
  rom[01729] = 16'h18c3;
  rom[01730] = 16'h10a2;
  rom[01731] = 16'h18a3;
  rom[01732] = 16'h10a2;
  rom[01733] = 16'h18c3;
  rom[01734] = 16'h10a2;
  rom[01735] = 16'h10a2;
  rom[01736] = 16'h10c2;
  rom[01737] = 16'h10a2;
  rom[01738] = 16'h18c3;
  rom[01739] = 16'h10a2;
  rom[01740] = 16'h18e3;
  rom[01741] = 16'hbdb6;
  rom[01742] = 16'hffdf;
  rom[01743] = 16'hffff;
  rom[01744] = 16'hffff;
  rom[01745] = 16'hffff;
  rom[01746] = 16'hffff;
  rom[01747] = 16'hffff;
  rom[01748] = 16'hffff;
  rom[01749] = 16'hffff;
  rom[01750] = 16'hffff;
  rom[01751] = 16'hffff;
  rom[01752] = 16'hffff;
  rom[01753] = 16'hffff;
  rom[01754] = 16'hffff;
  rom[01755] = 16'hffff;
  rom[01756] = 16'hffff;
  rom[01757] = 16'hffff;
  rom[01758] = 16'hffff;
  rom[01759] = 16'hffff;
  rom[01760] = 16'hffff;
  rom[01761] = 16'hffff;
  rom[01762] = 16'hffff;
  rom[01763] = 16'hffff;
  rom[01764] = 16'hffff;
  rom[01765] = 16'hffff;
  rom[01766] = 16'hffff;
  rom[01767] = 16'hffff;
  rom[01768] = 16'hffff;
  rom[01769] = 16'hffff;
  rom[01770] = 16'hffff;
  rom[01771] = 16'hffff;
  rom[01772] = 16'hffff;
  rom[01773] = 16'hffff;
  rom[01774] = 16'hffff;
  rom[01775] = 16'hffff;
  rom[01776] = 16'hffff;
  rom[01777] = 16'hffff;
  rom[01778] = 16'hffff;
  rom[01779] = 16'hffff;
  rom[01780] = 16'hffff;
  rom[01781] = 16'hffff;
  rom[01782] = 16'hffff;
  rom[01783] = 16'hffff;
  rom[01784] = 16'hffff;
  rom[01785] = 16'hffff;
  rom[01786] = 16'hffff;
  rom[01787] = 16'hffff;
  rom[01788] = 16'hffff;
  rom[01789] = 16'hffff;
  rom[01790] = 16'hffff;
  rom[01791] = 16'hffff;
  rom[01792] = 16'hffff;
  rom[01793] = 16'hffff;
  rom[01794] = 16'hffff;
  rom[01795] = 16'hffff;
  rom[01796] = 16'hffff;
  rom[01797] = 16'hffff;
  rom[01798] = 16'hffff;
  rom[01799] = 16'hffff;
  rom[01800] = 16'hffff;
  rom[01801] = 16'hffff;
  rom[01802] = 16'hffff;
  rom[01803] = 16'hffff;
  rom[01804] = 16'hffff;
  rom[01805] = 16'hffff;
  rom[01806] = 16'hffff;
  rom[01807] = 16'hffff;
  rom[01808] = 16'hffff;
  rom[01809] = 16'hffff;
  rom[01810] = 16'hffff;
  rom[01811] = 16'hffff;
  rom[01812] = 16'hffff;
  rom[01813] = 16'hffff;
  rom[01814] = 16'hffff;
  rom[01815] = 16'hffff;
  rom[01816] = 16'hffff;
  rom[01817] = 16'hffff;
  rom[01818] = 16'hffff;
  rom[01819] = 16'hffff;
  rom[01820] = 16'hffff;
  rom[01821] = 16'hffff;
  rom[01822] = 16'hffff;
  rom[01823] = 16'hffff;
  rom[01824] = 16'hffff;
  rom[01825] = 16'hffff;
  rom[01826] = 16'hffff;
  rom[01827] = 16'hffff;
  rom[01828] = 16'hffff;
  rom[01829] = 16'hffff;
  rom[01830] = 16'hffff;
  rom[01831] = 16'hffff;
  rom[01832] = 16'hffff;
  rom[01833] = 16'hffff;
  rom[01834] = 16'hffff;
  rom[01835] = 16'hffff;
  rom[01836] = 16'hffff;
  rom[01837] = 16'hffff;
  rom[01838] = 16'hffff;
  rom[01839] = 16'hffff;
  rom[01840] = 16'hffff;
  rom[01841] = 16'hffff;
  rom[01842] = 16'hffff;
  rom[01843] = 16'hffff;
  rom[01844] = 16'hffff;
  rom[01845] = 16'hffff;
  rom[01846] = 16'hffff;
  rom[01847] = 16'hffff;
  rom[01848] = 16'hffff;
  rom[01849] = 16'hffff;
  rom[01850] = 16'hffff;
  rom[01851] = 16'hffff;
  rom[01852] = 16'hffbe;
  rom[01853] = 16'h4a49;
  rom[01854] = 16'h18c2;
  rom[01855] = 16'h18c3;
  rom[01856] = 16'h18c3;
  rom[01857] = 16'h10a2;
  rom[01858] = 16'h18c3;
  rom[01859] = 16'h10a2;
  rom[01860] = 16'h18c3;
  rom[01861] = 16'h18a3;
  rom[01862] = 16'h18c3;
  rom[01863] = 16'h18c3;
  rom[01864] = 16'h18c3;
  rom[01865] = 16'h10c2;
  rom[01866] = 16'h18c3;
  rom[01867] = 16'h10a2;
  rom[01868] = 16'h18e3;
  rom[01869] = 16'h0861;
  rom[01870] = 16'h8c31;
  rom[01871] = 16'hffbe;
  rom[01872] = 16'hffff;
  rom[01873] = 16'hffff;
  rom[01874] = 16'hffff;
  rom[01875] = 16'hffff;
  rom[01876] = 16'hffff;
  rom[01877] = 16'hffff;
  rom[01878] = 16'hffff;
  rom[01879] = 16'hffff;
  rom[01880] = 16'hff9e;
  rom[01881] = 16'h734c;
  rom[01882] = 16'ha46f;
  rom[01883] = 16'h93eb;
  rom[01884] = 16'h8388;
  rom[01885] = 16'hde56;
  rom[01886] = 16'hffdf;
  rom[01887] = 16'hffdf;
  rom[01888] = 16'hffff;
  rom[01889] = 16'h9cd0;
  rom[01890] = 16'hc4cb;
  rom[01891] = 16'hf54a;
  rom[01892] = 16'hf56a;
  rom[01893] = 16'hfd49;
  rom[01894] = 16'hfd49;
  rom[01895] = 16'hfd48;
  rom[01896] = 16'hfd69;
  rom[01897] = 16'hfd48;
  rom[01898] = 16'hfd68;
  rom[01899] = 16'hf548;
  rom[01900] = 16'hfd48;
  rom[01901] = 16'hf548;
  rom[01902] = 16'hfd8b;
  rom[01903] = 16'hed6c;
  rom[01904] = 16'hc4cb;
  rom[01905] = 16'h6243;
  rom[01906] = 16'hde76;
  rom[01907] = 16'hd5d4;
  rom[01908] = 16'h9327;
  rom[01909] = 16'hdceb;
  rom[01910] = 16'he52b;
  rom[01911] = 16'hc4cc;
  rom[01912] = 16'h6266;
  rom[01913] = 16'hc5f5;
  rom[01914] = 16'hffff;
  rom[01915] = 16'hffff;
  rom[01916] = 16'hffff;
  rom[01917] = 16'hffdf;
  rom[01918] = 16'hdeba;
  rom[01919] = 16'hfffe;
  rom[01920] = 16'hfffe;
  rom[01921] = 16'hffff;
  rom[01922] = 16'hffbf;
  rom[01923] = 16'h83d0;
  rom[01924] = 16'h18e3;
  rom[01925] = 16'h10a2;
  rom[01926] = 16'h18a3;
  rom[01927] = 16'h10a2;
  rom[01928] = 16'h18c3;
  rom[01929] = 16'h10a2;
  rom[01930] = 16'h10a3;
  rom[01931] = 16'h10a2;
  rom[01932] = 16'h10a2;
  rom[01933] = 16'h10a2;
  rom[01934] = 16'h18c3;
  rom[01935] = 16'h10a2;
  rom[01936] = 16'h10c2;
  rom[01937] = 16'h18c2;
  rom[01938] = 16'h18c3;
  rom[01939] = 16'h10a2;
  rom[01940] = 16'h18a3;
  rom[01941] = 16'h8c51;
  rom[01942] = 16'hffbf;
  rom[01943] = 16'hffff;
  rom[01944] = 16'hffff;
  rom[01945] = 16'hffff;
  rom[01946] = 16'hffff;
  rom[01947] = 16'hffff;
  rom[01948] = 16'hffff;
  rom[01949] = 16'hffff;
  rom[01950] = 16'hffff;
  rom[01951] = 16'hffff;
  rom[01952] = 16'hffff;
  rom[01953] = 16'hffff;
  rom[01954] = 16'hffff;
  rom[01955] = 16'hffff;
  rom[01956] = 16'hffff;
  rom[01957] = 16'hffff;
  rom[01958] = 16'hffff;
  rom[01959] = 16'hffff;
  rom[01960] = 16'hffff;
  rom[01961] = 16'hffff;
  rom[01962] = 16'hffff;
  rom[01963] = 16'hffff;
  rom[01964] = 16'hffff;
  rom[01965] = 16'hffff;
  rom[01966] = 16'hffff;
  rom[01967] = 16'hffff;
  rom[01968] = 16'hffff;
  rom[01969] = 16'hffff;
  rom[01970] = 16'hffff;
  rom[01971] = 16'hffff;
  rom[01972] = 16'hffff;
  rom[01973] = 16'hffff;
  rom[01974] = 16'hffff;
  rom[01975] = 16'hffff;
  rom[01976] = 16'hffff;
  rom[01977] = 16'hffff;
  rom[01978] = 16'hffff;
  rom[01979] = 16'hffff;
  rom[01980] = 16'hffff;
  rom[01981] = 16'hffff;
  rom[01982] = 16'hffff;
  rom[01983] = 16'hffff;
  rom[01984] = 16'hffff;
  rom[01985] = 16'hffff;
  rom[01986] = 16'hffff;
  rom[01987] = 16'hffff;
  rom[01988] = 16'hffff;
  rom[01989] = 16'hffff;
  rom[01990] = 16'hffff;
  rom[01991] = 16'hffff;
  rom[01992] = 16'hffff;
  rom[01993] = 16'hffff;
  rom[01994] = 16'hffff;
  rom[01995] = 16'hffff;
  rom[01996] = 16'hffff;
  rom[01997] = 16'hffff;
  rom[01998] = 16'hffff;
  rom[01999] = 16'hffff;
  rom[02000] = 16'hffff;
  rom[02001] = 16'hffff;
  rom[02002] = 16'hffff;
  rom[02003] = 16'hffff;
  rom[02004] = 16'hffff;
  rom[02005] = 16'hffff;
  rom[02006] = 16'hffff;
  rom[02007] = 16'hffff;
  rom[02008] = 16'hffff;
  rom[02009] = 16'hffff;
  rom[02010] = 16'hffff;
  rom[02011] = 16'hffff;
  rom[02012] = 16'hffff;
  rom[02013] = 16'hffff;
  rom[02014] = 16'hffff;
  rom[02015] = 16'hffff;
  rom[02016] = 16'hffff;
  rom[02017] = 16'hffff;
  rom[02018] = 16'hffff;
  rom[02019] = 16'hffff;
  rom[02020] = 16'hffff;
  rom[02021] = 16'hffff;
  rom[02022] = 16'hffff;
  rom[02023] = 16'hffff;
  rom[02024] = 16'hffff;
  rom[02025] = 16'hffff;
  rom[02026] = 16'hffff;
  rom[02027] = 16'hffff;
  rom[02028] = 16'hffff;
  rom[02029] = 16'hffff;
  rom[02030] = 16'hffff;
  rom[02031] = 16'hffff;
  rom[02032] = 16'hffff;
  rom[02033] = 16'hffff;
  rom[02034] = 16'hffff;
  rom[02035] = 16'hffff;
  rom[02036] = 16'hffff;
  rom[02037] = 16'hffff;
  rom[02038] = 16'hffff;
  rom[02039] = 16'hffff;
  rom[02040] = 16'hffff;
  rom[02041] = 16'hffff;
  rom[02042] = 16'hffff;
  rom[02043] = 16'hffff;
  rom[02044] = 16'hffff;
  rom[02045] = 16'hffff;
  rom[02046] = 16'hffff;
  rom[02047] = 16'hffff;
  rom[02048] = 16'hffff;
  rom[02049] = 16'hffff;
  rom[02050] = 16'hffff;
  rom[02051] = 16'hffff;
  rom[02052] = 16'hdefb;
  rom[02053] = 16'h18e3;
  rom[02054] = 16'h0841;
  rom[02055] = 16'h20e4;
  rom[02056] = 16'h10a2;
  rom[02057] = 16'h10a2;
  rom[02058] = 16'h10a2;
  rom[02059] = 16'h10a2;
  rom[02060] = 16'h10a2;
  rom[02061] = 16'h18c3;
  rom[02062] = 16'h10a2;
  rom[02063] = 16'h10a2;
  rom[02064] = 16'h1082;
  rom[02065] = 16'h10c2;
  rom[02066] = 16'h10c2;
  rom[02067] = 16'h10a2;
  rom[02068] = 16'h10a2;
  rom[02069] = 16'h18c3;
  rom[02070] = 16'h6b6d;
  rom[02071] = 16'hffbf;
  rom[02072] = 16'hffff;
  rom[02073] = 16'hffff;
  rom[02074] = 16'hef5d;
  rom[02075] = 16'hdefb;
  rom[02076] = 16'hffff;
  rom[02077] = 16'hffff;
  rom[02078] = 16'hffff;
  rom[02079] = 16'hffff;
  rom[02080] = 16'hffdf;
  rom[02081] = 16'hb513;
  rom[02082] = 16'h7b29;
  rom[02083] = 16'hde12;
  rom[02084] = 16'h93e8;
  rom[02085] = 16'h9c2c;
  rom[02086] = 16'hf73b;
  rom[02087] = 16'hffff;
  rom[02088] = 16'hffdf;
  rom[02089] = 16'h9cb0;
  rom[02090] = 16'hc48a;
  rom[02091] = 16'hfd69;
  rom[02092] = 16'hf528;
  rom[02093] = 16'hfd68;
  rom[02094] = 16'hf548;
  rom[02095] = 16'hfd47;
  rom[02096] = 16'hf527;
  rom[02097] = 16'hfd68;
  rom[02098] = 16'hf548;
  rom[02099] = 16'hfd69;
  rom[02100] = 16'hfd69;
  rom[02101] = 16'hfd28;
  rom[02102] = 16'hf529;
  rom[02103] = 16'hf529;
  rom[02104] = 16'hdd4b;
  rom[02105] = 16'hac4a;
  rom[02106] = 16'h6aa5;
  rom[02107] = 16'h72c5;
  rom[02108] = 16'hbc08;
  rom[02109] = 16'hf52a;
  rom[02110] = 16'hed08;
  rom[02111] = 16'hf56d;
  rom[02112] = 16'hb46c;
  rom[02113] = 16'h8bec;
  rom[02114] = 16'hf77d;
  rom[02115] = 16'hffdf;
  rom[02116] = 16'hffdf;
  rom[02117] = 16'hf77d;
  rom[02118] = 16'h6b2a;
  rom[02119] = 16'h840d;
  rom[02120] = 16'he6f8;
  rom[02121] = 16'hfffe;
  rom[02122] = 16'hf77d;
  rom[02123] = 16'h7baf;
  rom[02124] = 16'h1082;
  rom[02125] = 16'h18c3;
  rom[02126] = 16'h10a3;
  rom[02127] = 16'h10a2;
  rom[02128] = 16'h10c2;
  rom[02129] = 16'h18e3;
  rom[02130] = 16'h10a2;
  rom[02131] = 16'h10c2;
  rom[02132] = 16'h10c2;
  rom[02133] = 16'h18c2;
  rom[02134] = 16'h10a2;
  rom[02135] = 16'h18c3;
  rom[02136] = 16'h18a2;
  rom[02137] = 16'h18e3;
  rom[02138] = 16'h0861;
  rom[02139] = 16'h18e3;
  rom[02140] = 16'h0861;
  rom[02141] = 16'h738e;
  rom[02142] = 16'hf77e;
  rom[02143] = 16'hffff;
  rom[02144] = 16'hffff;
  rom[02145] = 16'hffff;
  rom[02146] = 16'hffff;
  rom[02147] = 16'hffff;
  rom[02148] = 16'hffff;
  rom[02149] = 16'hffff;
  rom[02150] = 16'hffff;
  rom[02151] = 16'hffff;
  rom[02152] = 16'hffff;
  rom[02153] = 16'hffff;
  rom[02154] = 16'hffff;
  rom[02155] = 16'hffff;
  rom[02156] = 16'hffff;
  rom[02157] = 16'hffff;
  rom[02158] = 16'hffff;
  rom[02159] = 16'hffff;
  rom[02160] = 16'hffff;
  rom[02161] = 16'hffff;
  rom[02162] = 16'hffff;
  rom[02163] = 16'hffff;
  rom[02164] = 16'hffff;
  rom[02165] = 16'hffff;
  rom[02166] = 16'hffff;
  rom[02167] = 16'hffff;
  rom[02168] = 16'hffff;
  rom[02169] = 16'hffff;
  rom[02170] = 16'hffff;
  rom[02171] = 16'hffff;
  rom[02172] = 16'hffff;
  rom[02173] = 16'hffff;
  rom[02174] = 16'hffff;
  rom[02175] = 16'hffff;
  rom[02176] = 16'hffff;
  rom[02177] = 16'hffff;
  rom[02178] = 16'hffff;
  rom[02179] = 16'hffff;
  rom[02180] = 16'hffff;
  rom[02181] = 16'hffff;
  rom[02182] = 16'hffff;
  rom[02183] = 16'hffff;
  rom[02184] = 16'hffff;
  rom[02185] = 16'hffff;
  rom[02186] = 16'hffff;
  rom[02187] = 16'hffff;
  rom[02188] = 16'hffff;
  rom[02189] = 16'hffff;
  rom[02190] = 16'hffff;
  rom[02191] = 16'hffff;
  rom[02192] = 16'hffff;
  rom[02193] = 16'hffff;
  rom[02194] = 16'hffff;
  rom[02195] = 16'hffff;
  rom[02196] = 16'hffff;
  rom[02197] = 16'hffff;
  rom[02198] = 16'hffff;
  rom[02199] = 16'hffff;
  rom[02200] = 16'hffff;
  rom[02201] = 16'hffff;
  rom[02202] = 16'hffff;
  rom[02203] = 16'hffff;
  rom[02204] = 16'hffff;
  rom[02205] = 16'hffff;
  rom[02206] = 16'hffff;
  rom[02207] = 16'hffff;
  rom[02208] = 16'hffff;
  rom[02209] = 16'hffff;
  rom[02210] = 16'hffff;
  rom[02211] = 16'hffff;
  rom[02212] = 16'hffff;
  rom[02213] = 16'hffff;
  rom[02214] = 16'hffff;
  rom[02215] = 16'hffff;
  rom[02216] = 16'hffff;
  rom[02217] = 16'hffff;
  rom[02218] = 16'hffff;
  rom[02219] = 16'hffff;
  rom[02220] = 16'hffff;
  rom[02221] = 16'hffff;
  rom[02222] = 16'hffff;
  rom[02223] = 16'hffff;
  rom[02224] = 16'hffff;
  rom[02225] = 16'hffff;
  rom[02226] = 16'hffff;
  rom[02227] = 16'hffff;
  rom[02228] = 16'hffff;
  rom[02229] = 16'hffff;
  rom[02230] = 16'hffff;
  rom[02231] = 16'hffff;
  rom[02232] = 16'hffff;
  rom[02233] = 16'hffff;
  rom[02234] = 16'hffff;
  rom[02235] = 16'hffff;
  rom[02236] = 16'hffff;
  rom[02237] = 16'hffff;
  rom[02238] = 16'hffff;
  rom[02239] = 16'hffff;
  rom[02240] = 16'hffff;
  rom[02241] = 16'hffff;
  rom[02242] = 16'hffff;
  rom[02243] = 16'hffff;
  rom[02244] = 16'hffff;
  rom[02245] = 16'hffff;
  rom[02246] = 16'hffff;
  rom[02247] = 16'hffff;
  rom[02248] = 16'hffff;
  rom[02249] = 16'hffff;
  rom[02250] = 16'hffff;
  rom[02251] = 16'hffff;
  rom[02252] = 16'hce39;
  rom[02253] = 16'h10a2;
  rom[02254] = 16'h18c3;
  rom[02255] = 16'h0881;
  rom[02256] = 16'h18c3;
  rom[02257] = 16'h10a2;
  rom[02258] = 16'h18c3;
  rom[02259] = 16'h10a2;
  rom[02260] = 16'h18c3;
  rom[02261] = 16'h10a2;
  rom[02262] = 16'h18c3;
  rom[02263] = 16'h10a2;
  rom[02264] = 16'h18c3;
  rom[02265] = 16'h1082;
  rom[02266] = 16'h18c3;
  rom[02267] = 16'h10a2;
  rom[02268] = 16'h18c2;
  rom[02269] = 16'h10a2;
  rom[02270] = 16'h632d;
  rom[02271] = 16'hf77e;
  rom[02272] = 16'hffff;
  rom[02273] = 16'hffff;
  rom[02274] = 16'hce59;
  rom[02275] = 16'h73af;
  rom[02276] = 16'hef1c;
  rom[02277] = 16'hffff;
  rom[02278] = 16'hffff;
  rom[02279] = 16'hffff;
  rom[02280] = 16'hffff;
  rom[02281] = 16'hde98;
  rom[02282] = 16'h8b89;
  rom[02283] = 16'hcd4d;
  rom[02284] = 16'hd52d;
  rom[02285] = 16'h9368;
  rom[02286] = 16'hcdd5;
  rom[02287] = 16'hffdf;
  rom[02288] = 16'hffff;
  rom[02289] = 16'h942d;
  rom[02290] = 16'hccca;
  rom[02291] = 16'hfd6a;
  rom[02292] = 16'hfd49;
  rom[02293] = 16'hfd48;
  rom[02294] = 16'hfd68;
  rom[02295] = 16'hf547;
  rom[02296] = 16'hfd68;
  rom[02297] = 16'hfd47;
  rom[02298] = 16'hfd69;
  rom[02299] = 16'hfd48;
  rom[02300] = 16'hfd69;
  rom[02301] = 16'hfd48;
  rom[02302] = 16'hfd89;
  rom[02303] = 16'hf569;
  rom[02304] = 16'hed49;
  rom[02305] = 16'hedcd;
  rom[02306] = 16'hac08;
  rom[02307] = 16'hd4eb;
  rom[02308] = 16'hf54b;
  rom[02309] = 16'hfd28;
  rom[02310] = 16'hfd69;
  rom[02311] = 16'hed4a;
  rom[02312] = 16'hdd2e;
  rom[02313] = 16'h8b89;
  rom[02314] = 16'he678;
  rom[02315] = 16'hffdf;
  rom[02316] = 16'hffff;
  rom[02317] = 16'hdeb8;
  rom[02318] = 16'h6ae8;
  rom[02319] = 16'h940b;
  rom[02320] = 16'h8baa;
  rom[02321] = 16'hde35;
  rom[02322] = 16'hff9c;
  rom[02323] = 16'h7bce;
  rom[02324] = 16'h2124;
  rom[02325] = 16'h10c3;
  rom[02326] = 16'h10c2;
  rom[02327] = 16'h10c3;
  rom[02328] = 16'h18a3;
  rom[02329] = 16'h18c3;
  rom[02330] = 16'h18a3;
  rom[02331] = 16'h10a2;
  rom[02332] = 16'h10c3;
  rom[02333] = 16'h10a3;
  rom[02334] = 16'h18a3;
  rom[02335] = 16'h10a2;
  rom[02336] = 16'h18e3;
  rom[02337] = 16'h18c2;
  rom[02338] = 16'h1081;
  rom[02339] = 16'h10c2;
  rom[02340] = 16'h18c2;
  rom[02341] = 16'h6b4d;
  rom[02342] = 16'hffbf;
  rom[02343] = 16'hffff;
  rom[02344] = 16'hffff;
  rom[02345] = 16'hffff;
  rom[02346] = 16'hffff;
  rom[02347] = 16'hffff;
  rom[02348] = 16'hffff;
  rom[02349] = 16'hffff;
  rom[02350] = 16'hffff;
  rom[02351] = 16'hffff;
  rom[02352] = 16'hffff;
  rom[02353] = 16'hffff;
  rom[02354] = 16'hffff;
  rom[02355] = 16'hffff;
  rom[02356] = 16'hffff;
  rom[02357] = 16'hffff;
  rom[02358] = 16'hffff;
  rom[02359] = 16'hffff;
  rom[02360] = 16'hffff;
  rom[02361] = 16'hffff;
  rom[02362] = 16'hffff;
  rom[02363] = 16'hffff;
  rom[02364] = 16'hffff;
  rom[02365] = 16'hffff;
  rom[02366] = 16'hffff;
  rom[02367] = 16'hffff;
  rom[02368] = 16'hffff;
  rom[02369] = 16'hffff;
  rom[02370] = 16'hffff;
  rom[02371] = 16'hffff;
  rom[02372] = 16'hffff;
  rom[02373] = 16'hffff;
  rom[02374] = 16'hffff;
  rom[02375] = 16'hffff;
  rom[02376] = 16'hffff;
  rom[02377] = 16'hffff;
  rom[02378] = 16'hffff;
  rom[02379] = 16'hffff;
  rom[02380] = 16'hffff;
  rom[02381] = 16'hffff;
  rom[02382] = 16'hffff;
  rom[02383] = 16'hffff;
  rom[02384] = 16'hffff;
  rom[02385] = 16'hffff;
  rom[02386] = 16'hffff;
  rom[02387] = 16'hffff;
  rom[02388] = 16'hffff;
  rom[02389] = 16'hffff;
  rom[02390] = 16'hffff;
  rom[02391] = 16'hffff;
  rom[02392] = 16'hffff;
  rom[02393] = 16'hffff;
  rom[02394] = 16'hffff;
  rom[02395] = 16'hffff;
  rom[02396] = 16'hffff;
  rom[02397] = 16'hffff;
  rom[02398] = 16'hffff;
  rom[02399] = 16'hffff;
  rom[02400] = 16'hffff;
  rom[02401] = 16'hffff;
  rom[02402] = 16'hffff;
  rom[02403] = 16'hffff;
  rom[02404] = 16'hffff;
  rom[02405] = 16'hffff;
  rom[02406] = 16'hffff;
  rom[02407] = 16'hffff;
  rom[02408] = 16'hffff;
  rom[02409] = 16'hffff;
  rom[02410] = 16'hffff;
  rom[02411] = 16'hffff;
  rom[02412] = 16'hffff;
  rom[02413] = 16'hffff;
  rom[02414] = 16'hffff;
  rom[02415] = 16'hffff;
  rom[02416] = 16'hffff;
  rom[02417] = 16'hffff;
  rom[02418] = 16'hffff;
  rom[02419] = 16'hffff;
  rom[02420] = 16'hffff;
  rom[02421] = 16'hffff;
  rom[02422] = 16'hffff;
  rom[02423] = 16'hffff;
  rom[02424] = 16'hffff;
  rom[02425] = 16'hffff;
  rom[02426] = 16'hffff;
  rom[02427] = 16'hffff;
  rom[02428] = 16'hffff;
  rom[02429] = 16'hffff;
  rom[02430] = 16'hffff;
  rom[02431] = 16'hffff;
  rom[02432] = 16'hffff;
  rom[02433] = 16'hffff;
  rom[02434] = 16'hffff;
  rom[02435] = 16'hffff;
  rom[02436] = 16'hffff;
  rom[02437] = 16'hffff;
  rom[02438] = 16'hffff;
  rom[02439] = 16'hffff;
  rom[02440] = 16'hffff;
  rom[02441] = 16'hffff;
  rom[02442] = 16'hffff;
  rom[02443] = 16'hffff;
  rom[02444] = 16'hffff;
  rom[02445] = 16'hffff;
  rom[02446] = 16'hffff;
  rom[02447] = 16'hffff;
  rom[02448] = 16'hffff;
  rom[02449] = 16'hffff;
  rom[02450] = 16'hffff;
  rom[02451] = 16'hffff;
  rom[02452] = 16'hce38;
  rom[02453] = 16'h18a2;
  rom[02454] = 16'h18e3;
  rom[02455] = 16'h1081;
  rom[02456] = 16'h10a2;
  rom[02457] = 16'h10a2;
  rom[02458] = 16'h10a2;
  rom[02459] = 16'h10a2;
  rom[02460] = 16'h18c3;
  rom[02461] = 16'h10c2;
  rom[02462] = 16'h18c3;
  rom[02463] = 16'h10a2;
  rom[02464] = 16'h10c2;
  rom[02465] = 16'h18c3;
  rom[02466] = 16'h10a2;
  rom[02467] = 16'h10a2;
  rom[02468] = 16'h10c2;
  rom[02469] = 16'h10c3;
  rom[02470] = 16'h6b6e;
  rom[02471] = 16'hffbf;
  rom[02472] = 16'hfffe;
  rom[02473] = 16'hffff;
  rom[02474] = 16'he73d;
  rom[02475] = 16'h420a;
  rom[02476] = 16'h9491;
  rom[02477] = 16'hffde;
  rom[02478] = 16'hfffe;
  rom[02479] = 16'hffff;
  rom[02480] = 16'hfffe;
  rom[02481] = 16'hdeb8;
  rom[02482] = 16'h93e9;
  rom[02483] = 16'hc4ea;
  rom[02484] = 16'hedad;
  rom[02485] = 16'ha3c8;
  rom[02486] = 16'h93cb;
  rom[02487] = 16'hff5c;
  rom[02488] = 16'hffdd;
  rom[02489] = 16'h8b6a;
  rom[02490] = 16'hdcea;
  rom[02491] = 16'hfd6a;
  rom[02492] = 16'hfd48;
  rom[02493] = 16'hfd68;
  rom[02494] = 16'hfd48;
  rom[02495] = 16'hfd68;
  rom[02496] = 16'hf547;
  rom[02497] = 16'hfd67;
  rom[02498] = 16'hfd47;
  rom[02499] = 16'hfd68;
  rom[02500] = 16'hf548;
  rom[02501] = 16'hfd68;
  rom[02502] = 16'hfd88;
  rom[02503] = 16'hece5;
  rom[02504] = 16'hf5c9;
  rom[02505] = 16'hdca6;
  rom[02506] = 16'hf5cc;
  rom[02507] = 16'he50a;
  rom[02508] = 16'hf528;
  rom[02509] = 16'hfd69;
  rom[02510] = 16'hfd48;
  rom[02511] = 16'hf54a;
  rom[02512] = 16'he56d;
  rom[02513] = 16'h9bca;
  rom[02514] = 16'hddf6;
  rom[02515] = 16'hffff;
  rom[02516] = 16'hfffe;
  rom[02517] = 16'ha4cf;
  rom[02518] = 16'h93c9;
  rom[02519] = 16'hd590;
  rom[02520] = 16'ha3e9;
  rom[02521] = 16'h7b07;
  rom[02522] = 16'he676;
  rom[02523] = 16'ha4f2;
  rom[02524] = 16'h10e2;
  rom[02525] = 16'h10a2;
  rom[02526] = 16'h10c3;
  rom[02527] = 16'h10a2;
  rom[02528] = 16'h18e3;
  rom[02529] = 16'h1082;
  rom[02530] = 16'h18a3;
  rom[02531] = 16'h10a3;
  rom[02532] = 16'h10a3;
  rom[02533] = 16'h10a3;
  rom[02534] = 16'h18a3;
  rom[02535] = 16'h18a2;
  rom[02536] = 16'h10a2;
  rom[02537] = 16'h18a3;
  rom[02538] = 16'h1082;
  rom[02539] = 16'h18c3;
  rom[02540] = 16'h10a2;
  rom[02541] = 16'h6b4c;
  rom[02542] = 16'hf79e;
  rom[02543] = 16'hffff;
  rom[02544] = 16'hffff;
  rom[02545] = 16'hffff;
  rom[02546] = 16'hffff;
  rom[02547] = 16'hffff;
  rom[02548] = 16'hffff;
  rom[02549] = 16'hffff;
  rom[02550] = 16'hffff;
  rom[02551] = 16'hffff;
  rom[02552] = 16'hffff;
  rom[02553] = 16'hffff;
  rom[02554] = 16'hffff;
  rom[02555] = 16'hffff;
  rom[02556] = 16'hffff;
  rom[02557] = 16'hffff;
  rom[02558] = 16'hffff;
  rom[02559] = 16'hffff;
  rom[02560] = 16'hffff;
  rom[02561] = 16'hffff;
  rom[02562] = 16'hffff;
  rom[02563] = 16'hffff;
  rom[02564] = 16'hffff;
  rom[02565] = 16'hffff;
  rom[02566] = 16'hffff;
  rom[02567] = 16'hffff;
  rom[02568] = 16'hffff;
  rom[02569] = 16'hffff;
  rom[02570] = 16'hffff;
  rom[02571] = 16'hffff;
  rom[02572] = 16'hffff;
  rom[02573] = 16'hffff;
  rom[02574] = 16'hffff;
  rom[02575] = 16'hffff;
  rom[02576] = 16'hffff;
  rom[02577] = 16'hffff;
  rom[02578] = 16'hffff;
  rom[02579] = 16'hffff;
  rom[02580] = 16'hffff;
  rom[02581] = 16'hffff;
  rom[02582] = 16'hffff;
  rom[02583] = 16'hffff;
  rom[02584] = 16'hffff;
  rom[02585] = 16'hffff;
  rom[02586] = 16'hffff;
  rom[02587] = 16'hffff;
  rom[02588] = 16'hffff;
  rom[02589] = 16'hffff;
  rom[02590] = 16'hffff;
  rom[02591] = 16'hffff;
  rom[02592] = 16'hffff;
  rom[02593] = 16'hffff;
  rom[02594] = 16'hffff;
  rom[02595] = 16'hffff;
  rom[02596] = 16'hffff;
  rom[02597] = 16'hffff;
  rom[02598] = 16'hffff;
  rom[02599] = 16'hffff;
  rom[02600] = 16'hffff;
  rom[02601] = 16'hffff;
  rom[02602] = 16'hffff;
  rom[02603] = 16'hffff;
  rom[02604] = 16'hffff;
  rom[02605] = 16'hffff;
  rom[02606] = 16'hffff;
  rom[02607] = 16'hffff;
  rom[02608] = 16'hffff;
  rom[02609] = 16'hffff;
  rom[02610] = 16'hffff;
  rom[02611] = 16'hffff;
  rom[02612] = 16'hffff;
  rom[02613] = 16'hffff;
  rom[02614] = 16'hffff;
  rom[02615] = 16'hffff;
  rom[02616] = 16'hffff;
  rom[02617] = 16'hffff;
  rom[02618] = 16'hffff;
  rom[02619] = 16'hffff;
  rom[02620] = 16'hffff;
  rom[02621] = 16'hffff;
  rom[02622] = 16'hffff;
  rom[02623] = 16'hffff;
  rom[02624] = 16'hffff;
  rom[02625] = 16'hffff;
  rom[02626] = 16'hffff;
  rom[02627] = 16'hffff;
  rom[02628] = 16'hffff;
  rom[02629] = 16'hffff;
  rom[02630] = 16'hffff;
  rom[02631] = 16'hffff;
  rom[02632] = 16'hffff;
  rom[02633] = 16'hffff;
  rom[02634] = 16'hffff;
  rom[02635] = 16'hffff;
  rom[02636] = 16'hffff;
  rom[02637] = 16'hffff;
  rom[02638] = 16'hffff;
  rom[02639] = 16'hffff;
  rom[02640] = 16'hffff;
  rom[02641] = 16'hffff;
  rom[02642] = 16'hffff;
  rom[02643] = 16'hffff;
  rom[02644] = 16'hffff;
  rom[02645] = 16'hffff;
  rom[02646] = 16'hffff;
  rom[02647] = 16'hffff;
  rom[02648] = 16'hffff;
  rom[02649] = 16'hffff;
  rom[02650] = 16'hffff;
  rom[02651] = 16'hffff;
  rom[02652] = 16'hdeba;
  rom[02653] = 16'h10a1;
  rom[02654] = 16'h18c3;
  rom[02655] = 16'h18a2;
  rom[02656] = 16'h10a2;
  rom[02657] = 16'h1082;
  rom[02658] = 16'h18c3;
  rom[02659] = 16'h1082;
  rom[02660] = 16'h18c3;
  rom[02661] = 16'h10a2;
  rom[02662] = 16'h18c3;
  rom[02663] = 16'h18c3;
  rom[02664] = 16'h10a2;
  rom[02665] = 16'h10a2;
  rom[02666] = 16'h18a3;
  rom[02667] = 16'h18c3;
  rom[02668] = 16'h18c4;
  rom[02669] = 16'h10c3;
  rom[02670] = 16'h8411;
  rom[02671] = 16'hffbf;
  rom[02672] = 16'hffff;
  rom[02673] = 16'hffff;
  rom[02674] = 16'hf79f;
  rom[02675] = 16'h52ab;
  rom[02676] = 16'h4a08;
  rom[02677] = 16'hd658;
  rom[02678] = 16'hffff;
  rom[02679] = 16'hffff;
  rom[02680] = 16'hffff;
  rom[02681] = 16'he6f9;
  rom[02682] = 16'h9bea;
  rom[02683] = 16'hdd6b;
  rom[02684] = 16'hed6a;
  rom[02685] = 16'hd50b;
  rom[02686] = 16'h7a85;
  rom[02687] = 16'he677;
  rom[02688] = 16'hde57;
  rom[02689] = 16'h8307;
  rom[02690] = 16'he52b;
  rom[02691] = 16'hfd69;
  rom[02692] = 16'hfd69;
  rom[02693] = 16'hfd68;
  rom[02694] = 16'hfd68;
  rom[02695] = 16'hfd68;
  rom[02696] = 16'hfd68;
  rom[02697] = 16'hfd67;
  rom[02698] = 16'hfd68;
  rom[02699] = 16'hfd68;
  rom[02700] = 16'hfd69;
  rom[02701] = 16'hfd48;
  rom[02702] = 16'hfd69;
  rom[02703] = 16'hfd88;
  rom[02704] = 16'hf568;
  rom[02705] = 16'hf589;
  rom[02706] = 16'hf56a;
  rom[02707] = 16'hfdcb;
  rom[02708] = 16'hfd69;
  rom[02709] = 16'hf547;
  rom[02710] = 16'hfd48;
  rom[02711] = 16'hf54a;
  rom[02712] = 16'hedae;
  rom[02713] = 16'h9bc8;
  rom[02714] = 16'hc511;
  rom[02715] = 16'hffde;
  rom[02716] = 16'hf71a;
  rom[02717] = 16'h6a64;
  rom[02718] = 16'hc4ac;
  rom[02719] = 16'hed8e;
  rom[02720] = 16'he56e;
  rom[02721] = 16'ha3c8;
  rom[02722] = 16'h8348;
  rom[02723] = 16'ha4b0;
  rom[02724] = 16'h18c2;
  rom[02725] = 16'h10c3;
  rom[02726] = 16'h10e3;
  rom[02727] = 16'h08a2;
  rom[02728] = 16'h18c3;
  rom[02729] = 16'h18a2;
  rom[02730] = 16'h18a3;
  rom[02731] = 16'h10a2;
  rom[02732] = 16'h10c2;
  rom[02733] = 16'h10c2;
  rom[02734] = 16'h18a2;
  rom[02735] = 16'h18a2;
  rom[02736] = 16'h18a3;
  rom[02737] = 16'h18a2;
  rom[02738] = 16'h1082;
  rom[02739] = 16'h18c3;
  rom[02740] = 16'h18c2;
  rom[02741] = 16'h7bcf;
  rom[02742] = 16'hffbf;
  rom[02743] = 16'hffff;
  rom[02744] = 16'hffff;
  rom[02745] = 16'hffff;
  rom[02746] = 16'hffff;
  rom[02747] = 16'hffff;
  rom[02748] = 16'hffff;
  rom[02749] = 16'hffff;
  rom[02750] = 16'hffff;
  rom[02751] = 16'hffff;
  rom[02752] = 16'hffff;
  rom[02753] = 16'hffff;
  rom[02754] = 16'hffff;
  rom[02755] = 16'hffff;
  rom[02756] = 16'hffff;
  rom[02757] = 16'hffff;
  rom[02758] = 16'hffff;
  rom[02759] = 16'hffff;
  rom[02760] = 16'hffff;
  rom[02761] = 16'hffff;
  rom[02762] = 16'hffff;
  rom[02763] = 16'hffff;
  rom[02764] = 16'hffff;
  rom[02765] = 16'hffff;
  rom[02766] = 16'hffff;
  rom[02767] = 16'hffff;
  rom[02768] = 16'hffff;
  rom[02769] = 16'hffff;
  rom[02770] = 16'hffff;
  rom[02771] = 16'hffff;
  rom[02772] = 16'hffff;
  rom[02773] = 16'hffff;
  rom[02774] = 16'hffff;
  rom[02775] = 16'hffff;
  rom[02776] = 16'hffff;
  rom[02777] = 16'hffff;
  rom[02778] = 16'hffff;
  rom[02779] = 16'hffff;
  rom[02780] = 16'hffff;
  rom[02781] = 16'hffff;
  rom[02782] = 16'hffff;
  rom[02783] = 16'hffff;
  rom[02784] = 16'hffff;
  rom[02785] = 16'hffff;
  rom[02786] = 16'hffff;
  rom[02787] = 16'hffff;
  rom[02788] = 16'hffff;
  rom[02789] = 16'hffff;
  rom[02790] = 16'hffff;
  rom[02791] = 16'hffff;
  rom[02792] = 16'hffff;
  rom[02793] = 16'hffff;
  rom[02794] = 16'hffff;
  rom[02795] = 16'hffff;
  rom[02796] = 16'hffff;
  rom[02797] = 16'hffff;
  rom[02798] = 16'hffff;
  rom[02799] = 16'hffff;
  rom[02800] = 16'hffff;
  rom[02801] = 16'hffff;
  rom[02802] = 16'hffff;
  rom[02803] = 16'hffff;
  rom[02804] = 16'hffff;
  rom[02805] = 16'hffff;
  rom[02806] = 16'hffff;
  rom[02807] = 16'hffff;
  rom[02808] = 16'hffff;
  rom[02809] = 16'hffff;
  rom[02810] = 16'hffff;
  rom[02811] = 16'hffff;
  rom[02812] = 16'hffff;
  rom[02813] = 16'hffff;
  rom[02814] = 16'hffff;
  rom[02815] = 16'hffff;
  rom[02816] = 16'hffff;
  rom[02817] = 16'hffff;
  rom[02818] = 16'hffff;
  rom[02819] = 16'hffff;
  rom[02820] = 16'hffff;
  rom[02821] = 16'hffff;
  rom[02822] = 16'hffff;
  rom[02823] = 16'hffff;
  rom[02824] = 16'hffff;
  rom[02825] = 16'hffff;
  rom[02826] = 16'hffff;
  rom[02827] = 16'hffff;
  rom[02828] = 16'hffff;
  rom[02829] = 16'hffff;
  rom[02830] = 16'hffff;
  rom[02831] = 16'hffff;
  rom[02832] = 16'hffff;
  rom[02833] = 16'hffff;
  rom[02834] = 16'hffff;
  rom[02835] = 16'hffff;
  rom[02836] = 16'hffff;
  rom[02837] = 16'hffff;
  rom[02838] = 16'hffff;
  rom[02839] = 16'hffff;
  rom[02840] = 16'hffff;
  rom[02841] = 16'hffff;
  rom[02842] = 16'hffff;
  rom[02843] = 16'hffff;
  rom[02844] = 16'hffff;
  rom[02845] = 16'hffff;
  rom[02846] = 16'hffff;
  rom[02847] = 16'hffff;
  rom[02848] = 16'hffff;
  rom[02849] = 16'hffff;
  rom[02850] = 16'hffff;
  rom[02851] = 16'hffff;
  rom[02852] = 16'hef5d;
  rom[02853] = 16'h3165;
  rom[02854] = 16'h1082;
  rom[02855] = 16'h18e3;
  rom[02856] = 16'h10a2;
  rom[02857] = 16'h1082;
  rom[02858] = 16'h10a2;
  rom[02859] = 16'h10a2;
  rom[02860] = 16'h10a2;
  rom[02861] = 16'h18c3;
  rom[02862] = 16'h10a2;
  rom[02863] = 16'h18c3;
  rom[02864] = 16'h0861;
  rom[02865] = 16'h10c2;
  rom[02866] = 16'h10a2;
  rom[02867] = 16'h10a2;
  rom[02868] = 16'h1083;
  rom[02869] = 16'h0882;
  rom[02870] = 16'h9492;
  rom[02871] = 16'hff9f;
  rom[02872] = 16'hffde;
  rom[02873] = 16'hffff;
  rom[02874] = 16'hf7be;
  rom[02875] = 16'h8c30;
  rom[02876] = 16'h83ac;
  rom[02877] = 16'h83ae;
  rom[02878] = 16'hff7e;
  rom[02879] = 16'hffbf;
  rom[02880] = 16'hf77e;
  rom[02881] = 16'hf71a;
  rom[02882] = 16'h93a9;
  rom[02883] = 16'hdd4a;
  rom[02884] = 16'hed88;
  rom[02885] = 16'hed8a;
  rom[02886] = 16'ha386;
  rom[02887] = 16'h59e3;
  rom[02888] = 16'h61e3;
  rom[02889] = 16'habe8;
  rom[02890] = 16'hed4a;
  rom[02891] = 16'hf548;
  rom[02892] = 16'hf548;
  rom[02893] = 16'hfd68;
  rom[02894] = 16'hf547;
  rom[02895] = 16'hf568;
  rom[02896] = 16'hfd68;
  rom[02897] = 16'hfd88;
  rom[02898] = 16'hf568;
  rom[02899] = 16'hfd88;
  rom[02900] = 16'hfd68;
  rom[02901] = 16'hfd49;
  rom[02902] = 16'hfd29;
  rom[02903] = 16'hf527;
  rom[02904] = 16'hfd88;
  rom[02905] = 16'hf547;
  rom[02906] = 16'hed68;
  rom[02907] = 16'hf568;
  rom[02908] = 16'hf527;
  rom[02909] = 16'hfda8;
  rom[02910] = 16'hed27;
  rom[02911] = 16'hf58b;
  rom[02912] = 16'he56c;
  rom[02913] = 16'h9bc7;
  rom[02914] = 16'hac8d;
  rom[02915] = 16'hf719;
  rom[02916] = 16'h82e8;
  rom[02917] = 16'h9305;
  rom[02918] = 16'hed6d;
  rom[02919] = 16'he4ea;
  rom[02920] = 16'hed4b;
  rom[02921] = 16'he52c;
  rom[02922] = 16'ha3e8;
  rom[02923] = 16'h72c8;
  rom[02924] = 16'h5208;
  rom[02925] = 16'h1062;
  rom[02926] = 16'h10c2;
  rom[02927] = 16'h10c3;
  rom[02928] = 16'h1082;
  rom[02929] = 16'h18a3;
  rom[02930] = 16'h18a2;
  rom[02931] = 16'h10a2;
  rom[02932] = 16'h10c2;
  rom[02933] = 16'h10c2;
  rom[02934] = 16'h18a2;
  rom[02935] = 16'h1081;
  rom[02936] = 16'h18a3;
  rom[02937] = 16'h10a2;
  rom[02938] = 16'h10a1;
  rom[02939] = 16'h10a2;
  rom[02940] = 16'h0861;
  rom[02941] = 16'h9cf3;
  rom[02942] = 16'hffdf;
  rom[02943] = 16'hffff;
  rom[02944] = 16'hffff;
  rom[02945] = 16'hffff;
  rom[02946] = 16'hffff;
  rom[02947] = 16'hffff;
  rom[02948] = 16'hffff;
  rom[02949] = 16'hffff;
  rom[02950] = 16'hffff;
  rom[02951] = 16'hffff;
  rom[02952] = 16'hffff;
  rom[02953] = 16'hffff;
  rom[02954] = 16'hffff;
  rom[02955] = 16'hffff;
  rom[02956] = 16'hffff;
  rom[02957] = 16'hffff;
  rom[02958] = 16'hffff;
  rom[02959] = 16'hffff;
  rom[02960] = 16'hffff;
  rom[02961] = 16'hffff;
  rom[02962] = 16'hffff;
  rom[02963] = 16'hffff;
  rom[02964] = 16'hffff;
  rom[02965] = 16'hffff;
  rom[02966] = 16'hffff;
  rom[02967] = 16'hffff;
  rom[02968] = 16'hffff;
  rom[02969] = 16'hffff;
  rom[02970] = 16'hffff;
  rom[02971] = 16'hffff;
  rom[02972] = 16'hffff;
  rom[02973] = 16'hffff;
  rom[02974] = 16'hffff;
  rom[02975] = 16'hffff;
  rom[02976] = 16'hffff;
  rom[02977] = 16'hffff;
  rom[02978] = 16'hffff;
  rom[02979] = 16'hffff;
  rom[02980] = 16'hffff;
  rom[02981] = 16'hffff;
  rom[02982] = 16'hffff;
  rom[02983] = 16'hffff;
  rom[02984] = 16'hffff;
  rom[02985] = 16'hffff;
  rom[02986] = 16'hffff;
  rom[02987] = 16'hffff;
  rom[02988] = 16'hffff;
  rom[02989] = 16'hffff;
  rom[02990] = 16'hffff;
  rom[02991] = 16'hffff;
  rom[02992] = 16'hffff;
  rom[02993] = 16'hffff;
  rom[02994] = 16'hffff;
  rom[02995] = 16'hffff;
  rom[02996] = 16'hffff;
  rom[02997] = 16'hffff;
  rom[02998] = 16'hffff;
  rom[02999] = 16'hffff;
  rom[03000] = 16'hffff;
  rom[03001] = 16'hffff;
  rom[03002] = 16'hffff;
  rom[03003] = 16'hffff;
  rom[03004] = 16'hffff;
  rom[03005] = 16'hffff;
  rom[03006] = 16'hffff;
  rom[03007] = 16'hffff;
  rom[03008] = 16'hffff;
  rom[03009] = 16'hffff;
  rom[03010] = 16'hffff;
  rom[03011] = 16'hffff;
  rom[03012] = 16'hffff;
  rom[03013] = 16'hffff;
  rom[03014] = 16'hffff;
  rom[03015] = 16'hffff;
  rom[03016] = 16'hffff;
  rom[03017] = 16'hffff;
  rom[03018] = 16'hffff;
  rom[03019] = 16'hffff;
  rom[03020] = 16'hffff;
  rom[03021] = 16'hffff;
  rom[03022] = 16'hffff;
  rom[03023] = 16'hffff;
  rom[03024] = 16'hffff;
  rom[03025] = 16'hffff;
  rom[03026] = 16'hffff;
  rom[03027] = 16'hffff;
  rom[03028] = 16'hffff;
  rom[03029] = 16'hffff;
  rom[03030] = 16'hffff;
  rom[03031] = 16'hffff;
  rom[03032] = 16'hffff;
  rom[03033] = 16'hffff;
  rom[03034] = 16'hffff;
  rom[03035] = 16'hffff;
  rom[03036] = 16'hffff;
  rom[03037] = 16'hffff;
  rom[03038] = 16'hffff;
  rom[03039] = 16'hffff;
  rom[03040] = 16'hffff;
  rom[03041] = 16'hffff;
  rom[03042] = 16'hffff;
  rom[03043] = 16'hffff;
  rom[03044] = 16'hffff;
  rom[03045] = 16'hffff;
  rom[03046] = 16'hffff;
  rom[03047] = 16'hffff;
  rom[03048] = 16'hffff;
  rom[03049] = 16'hffff;
  rom[03050] = 16'hffff;
  rom[03051] = 16'hffff;
  rom[03052] = 16'hffdf;
  rom[03053] = 16'h62ec;
  rom[03054] = 16'h1082;
  rom[03055] = 16'h18e2;
  rom[03056] = 16'h18e3;
  rom[03057] = 16'h1082;
  rom[03058] = 16'h18c3;
  rom[03059] = 16'h18c3;
  rom[03060] = 16'h10a2;
  rom[03061] = 16'h18a3;
  rom[03062] = 16'h18c3;
  rom[03063] = 16'h10a2;
  rom[03064] = 16'h18e3;
  rom[03065] = 16'h18a3;
  rom[03066] = 16'h10a2;
  rom[03067] = 16'h10a2;
  rom[03068] = 16'h18c3;
  rom[03069] = 16'h2144;
  rom[03070] = 16'hbdf7;
  rom[03071] = 16'hffff;
  rom[03072] = 16'hffff;
  rom[03073] = 16'hffde;
  rom[03074] = 16'hfffe;
  rom[03075] = 16'h9caf;
  rom[03076] = 16'hbd31;
  rom[03077] = 16'h6aa8;
  rom[03078] = 16'he69b;
  rom[03079] = 16'hf75e;
  rom[03080] = 16'hffff;
  rom[03081] = 16'hc553;
  rom[03082] = 16'h9347;
  rom[03083] = 16'he529;
  rom[03084] = 16'hfda8;
  rom[03085] = 16'hf569;
  rom[03086] = 16'he54b;
  rom[03087] = 16'hccab;
  rom[03088] = 16'hdd2d;
  rom[03089] = 16'he54c;
  rom[03090] = 16'hfdab;
  rom[03091] = 16'hf568;
  rom[03092] = 16'hfda9;
  rom[03093] = 16'hfd68;
  rom[03094] = 16'hfd89;
  rom[03095] = 16'hfd88;
  rom[03096] = 16'hfd89;
  rom[03097] = 16'hfd68;
  rom[03098] = 16'hfd89;
  rom[03099] = 16'hfd68;
  rom[03100] = 16'hfd89;
  rom[03101] = 16'hfd48;
  rom[03102] = 16'hfd6a;
  rom[03103] = 16'hfd68;
  rom[03104] = 16'hfd27;
  rom[03105] = 16'hfd87;
  rom[03106] = 16'hfd88;
  rom[03107] = 16'hfd68;
  rom[03108] = 16'hfd88;
  rom[03109] = 16'hfd87;
  rom[03110] = 16'hf568;
  rom[03111] = 16'hf58a;
  rom[03112] = 16'he56b;
  rom[03113] = 16'hbc68;
  rom[03114] = 16'h82a4;
  rom[03115] = 16'h69e3;
  rom[03116] = 16'ha388;
  rom[03117] = 16'hed6d;
  rom[03118] = 16'hf50a;
  rom[03119] = 16'hf549;
  rom[03120] = 16'hfd29;
  rom[03121] = 16'hed6a;
  rom[03122] = 16'he54d;
  rom[03123] = 16'h82e6;
  rom[03124] = 16'h51c5;
  rom[03125] = 16'h20c2;
  rom[03126] = 16'h1082;
  rom[03127] = 16'h10a3;
  rom[03128] = 16'h18c3;
  rom[03129] = 16'h18a3;
  rom[03130] = 16'h18a2;
  rom[03131] = 16'h10a2;
  rom[03132] = 16'h10c2;
  rom[03133] = 16'h10c2;
  rom[03134] = 16'h18a2;
  rom[03135] = 16'h18c2;
  rom[03136] = 16'h18a2;
  rom[03137] = 16'h1082;
  rom[03138] = 16'h2124;
  rom[03139] = 16'h10a2;
  rom[03140] = 16'h2945;
  rom[03141] = 16'hc618;
  rom[03142] = 16'hffff;
  rom[03143] = 16'hffff;
  rom[03144] = 16'hffff;
  rom[03145] = 16'hffff;
  rom[03146] = 16'hffff;
  rom[03147] = 16'hffff;
  rom[03148] = 16'hffff;
  rom[03149] = 16'hffff;
  rom[03150] = 16'hffff;
  rom[03151] = 16'hffff;
  rom[03152] = 16'hffff;
  rom[03153] = 16'hffff;
  rom[03154] = 16'hffff;
  rom[03155] = 16'hffff;
  rom[03156] = 16'hffff;
  rom[03157] = 16'hffff;
  rom[03158] = 16'hffff;
  rom[03159] = 16'hffff;
  rom[03160] = 16'hffff;
  rom[03161] = 16'hffff;
  rom[03162] = 16'hffff;
  rom[03163] = 16'hffff;
  rom[03164] = 16'hffff;
  rom[03165] = 16'hffff;
  rom[03166] = 16'hffff;
  rom[03167] = 16'hffff;
  rom[03168] = 16'hffff;
  rom[03169] = 16'hffff;
  rom[03170] = 16'hffff;
  rom[03171] = 16'hffff;
  rom[03172] = 16'hffff;
  rom[03173] = 16'hffff;
  rom[03174] = 16'hffff;
  rom[03175] = 16'hffff;
  rom[03176] = 16'hffff;
  rom[03177] = 16'hffff;
  rom[03178] = 16'hffff;
  rom[03179] = 16'hffff;
  rom[03180] = 16'hffff;
  rom[03181] = 16'hffff;
  rom[03182] = 16'hffff;
  rom[03183] = 16'hffff;
  rom[03184] = 16'hffff;
  rom[03185] = 16'hffff;
  rom[03186] = 16'hffff;
  rom[03187] = 16'hffff;
  rom[03188] = 16'hffff;
  rom[03189] = 16'hffff;
  rom[03190] = 16'hffff;
  rom[03191] = 16'hffff;
  rom[03192] = 16'hffff;
  rom[03193] = 16'hffff;
  rom[03194] = 16'hffff;
  rom[03195] = 16'hffff;
  rom[03196] = 16'hffff;
  rom[03197] = 16'hffff;
  rom[03198] = 16'hffff;
  rom[03199] = 16'hffff;
  rom[03200] = 16'hffff;
  rom[03201] = 16'hffff;
  rom[03202] = 16'hffff;
  rom[03203] = 16'hffff;
  rom[03204] = 16'hffff;
  rom[03205] = 16'hffff;
  rom[03206] = 16'hffff;
  rom[03207] = 16'hffff;
  rom[03208] = 16'hffff;
  rom[03209] = 16'hffff;
  rom[03210] = 16'hffff;
  rom[03211] = 16'hffff;
  rom[03212] = 16'hffff;
  rom[03213] = 16'hffff;
  rom[03214] = 16'hffff;
  rom[03215] = 16'hffff;
  rom[03216] = 16'hffff;
  rom[03217] = 16'hffff;
  rom[03218] = 16'hffff;
  rom[03219] = 16'hffff;
  rom[03220] = 16'hffff;
  rom[03221] = 16'hffff;
  rom[03222] = 16'hffff;
  rom[03223] = 16'hffff;
  rom[03224] = 16'hffff;
  rom[03225] = 16'hffff;
  rom[03226] = 16'hffff;
  rom[03227] = 16'hffff;
  rom[03228] = 16'hffff;
  rom[03229] = 16'hffff;
  rom[03230] = 16'hffff;
  rom[03231] = 16'hffff;
  rom[03232] = 16'hffff;
  rom[03233] = 16'hffff;
  rom[03234] = 16'hffff;
  rom[03235] = 16'hffff;
  rom[03236] = 16'hffff;
  rom[03237] = 16'hffff;
  rom[03238] = 16'hffff;
  rom[03239] = 16'hffff;
  rom[03240] = 16'hffff;
  rom[03241] = 16'hffff;
  rom[03242] = 16'hffff;
  rom[03243] = 16'hffff;
  rom[03244] = 16'hffff;
  rom[03245] = 16'hffff;
  rom[03246] = 16'hffff;
  rom[03247] = 16'hffff;
  rom[03248] = 16'hffff;
  rom[03249] = 16'hffff;
  rom[03250] = 16'hffff;
  rom[03251] = 16'hffff;
  rom[03252] = 16'hffde;
  rom[03253] = 16'ha4f4;
  rom[03254] = 16'h18c2;
  rom[03255] = 16'h1082;
  rom[03256] = 16'h10c2;
  rom[03257] = 16'h10a2;
  rom[03258] = 16'h10a2;
  rom[03259] = 16'h10a2;
  rom[03260] = 16'h10a2;
  rom[03261] = 16'h10a2;
  rom[03262] = 16'h10a2;
  rom[03263] = 16'h18a3;
  rom[03264] = 16'h10c2;
  rom[03265] = 16'h10a2;
  rom[03266] = 16'h18c3;
  rom[03267] = 16'h18c3;
  rom[03268] = 16'h10a2;
  rom[03269] = 16'h52ea;
  rom[03270] = 16'he75b;
  rom[03271] = 16'hffff;
  rom[03272] = 16'hffde;
  rom[03273] = 16'hfffe;
  rom[03274] = 16'hffdd;
  rom[03275] = 16'h9cad;
  rom[03276] = 16'haccc;
  rom[03277] = 16'h9c0b;
  rom[03278] = 16'ha470;
  rom[03279] = 16'hffdf;
  rom[03280] = 16'hf73a;
  rom[03281] = 16'h7b07;
  rom[03282] = 16'hb449;
  rom[03283] = 16'hf58b;
  rom[03284] = 16'hf547;
  rom[03285] = 16'hfd68;
  rom[03286] = 16'hfd8a;
  rom[03287] = 16'hed4b;
  rom[03288] = 16'hed6b;
  rom[03289] = 16'hf56a;
  rom[03290] = 16'hfda9;
  rom[03291] = 16'hf568;
  rom[03292] = 16'hf588;
  rom[03293] = 16'hfd68;
  rom[03294] = 16'hfd68;
  rom[03295] = 16'hfd88;
  rom[03296] = 16'hf568;
  rom[03297] = 16'hfd88;
  rom[03298] = 16'hfd68;
  rom[03299] = 16'hfd88;
  rom[03300] = 16'hf568;
  rom[03301] = 16'hfd69;
  rom[03302] = 16'hfd68;
  rom[03303] = 16'hfd68;
  rom[03304] = 16'hf567;
  rom[03305] = 16'hfd88;
  rom[03306] = 16'hfd47;
  rom[03307] = 16'hfd47;
  rom[03308] = 16'hfd67;
  rom[03309] = 16'hfd67;
  rom[03310] = 16'hf547;
  rom[03311] = 16'hf569;
  rom[03312] = 16'hed6a;
  rom[03313] = 16'hedab;
  rom[03314] = 16'hd4eb;
  rom[03315] = 16'hed6d;
  rom[03316] = 16'hed4b;
  rom[03317] = 16'hf56a;
  rom[03318] = 16'hfd69;
  rom[03319] = 16'hfd28;
  rom[03320] = 16'hf527;
  rom[03321] = 16'hfd8a;
  rom[03322] = 16'he52b;
  rom[03323] = 16'hcced;
  rom[03324] = 16'h51c3;
  rom[03325] = 16'h30e1;
  rom[03326] = 16'h1881;
  rom[03327] = 16'h18c3;
  rom[03328] = 16'h10a3;
  rom[03329] = 16'h18a3;
  rom[03330] = 16'h1882;
  rom[03331] = 16'h10a2;
  rom[03332] = 16'h10a2;
  rom[03333] = 16'h10c2;
  rom[03334] = 16'h18a2;
  rom[03335] = 16'h18c2;
  rom[03336] = 16'h10a2;
  rom[03337] = 16'h18c2;
  rom[03338] = 16'h10a2;
  rom[03339] = 16'h18c3;
  rom[03340] = 16'h5aeb;
  rom[03341] = 16'hf75e;
  rom[03342] = 16'hffff;
  rom[03343] = 16'hffff;
  rom[03344] = 16'hffff;
  rom[03345] = 16'hffff;
  rom[03346] = 16'hffff;
  rom[03347] = 16'hffff;
  rom[03348] = 16'hffff;
  rom[03349] = 16'hffff;
  rom[03350] = 16'hffff;
  rom[03351] = 16'hffff;
  rom[03352] = 16'hffff;
  rom[03353] = 16'hffff;
  rom[03354] = 16'hffff;
  rom[03355] = 16'hffff;
  rom[03356] = 16'hffff;
  rom[03357] = 16'hffff;
  rom[03358] = 16'hffff;
  rom[03359] = 16'hffff;
  rom[03360] = 16'hffff;
  rom[03361] = 16'hffff;
  rom[03362] = 16'hffff;
  rom[03363] = 16'hffff;
  rom[03364] = 16'hffff;
  rom[03365] = 16'hffff;
  rom[03366] = 16'hffff;
  rom[03367] = 16'hffff;
  rom[03368] = 16'hffff;
  rom[03369] = 16'hffff;
  rom[03370] = 16'hffff;
  rom[03371] = 16'hffff;
  rom[03372] = 16'hffff;
  rom[03373] = 16'hffff;
  rom[03374] = 16'hffff;
  rom[03375] = 16'hffff;
  rom[03376] = 16'hffff;
  rom[03377] = 16'hffff;
  rom[03378] = 16'hffff;
  rom[03379] = 16'hffff;
  rom[03380] = 16'hffff;
  rom[03381] = 16'hffff;
  rom[03382] = 16'hffff;
  rom[03383] = 16'hffff;
  rom[03384] = 16'hffff;
  rom[03385] = 16'hffff;
  rom[03386] = 16'hffff;
  rom[03387] = 16'hffff;
  rom[03388] = 16'hffff;
  rom[03389] = 16'hffff;
  rom[03390] = 16'hffff;
  rom[03391] = 16'hffff;
  rom[03392] = 16'hffff;
  rom[03393] = 16'hffff;
  rom[03394] = 16'hffff;
  rom[03395] = 16'hffff;
  rom[03396] = 16'hffff;
  rom[03397] = 16'hffff;
  rom[03398] = 16'hffff;
  rom[03399] = 16'hffff;
  rom[03400] = 16'hffff;
  rom[03401] = 16'hffff;
  rom[03402] = 16'hffff;
  rom[03403] = 16'hffff;
  rom[03404] = 16'hffff;
  rom[03405] = 16'hffff;
  rom[03406] = 16'hffff;
  rom[03407] = 16'hffff;
  rom[03408] = 16'hffff;
  rom[03409] = 16'hffff;
  rom[03410] = 16'hffff;
  rom[03411] = 16'hffff;
  rom[03412] = 16'hffff;
  rom[03413] = 16'hffff;
  rom[03414] = 16'hffff;
  rom[03415] = 16'hffff;
  rom[03416] = 16'hffff;
  rom[03417] = 16'hffff;
  rom[03418] = 16'hffff;
  rom[03419] = 16'hffff;
  rom[03420] = 16'hffff;
  rom[03421] = 16'hffff;
  rom[03422] = 16'hffff;
  rom[03423] = 16'hffff;
  rom[03424] = 16'hffff;
  rom[03425] = 16'hffff;
  rom[03426] = 16'hffff;
  rom[03427] = 16'hffff;
  rom[03428] = 16'hffff;
  rom[03429] = 16'hffff;
  rom[03430] = 16'hffff;
  rom[03431] = 16'hffff;
  rom[03432] = 16'hffff;
  rom[03433] = 16'hffff;
  rom[03434] = 16'hffff;
  rom[03435] = 16'hffff;
  rom[03436] = 16'hffff;
  rom[03437] = 16'hffff;
  rom[03438] = 16'hffff;
  rom[03439] = 16'hffff;
  rom[03440] = 16'hffff;
  rom[03441] = 16'hffff;
  rom[03442] = 16'hffff;
  rom[03443] = 16'hffff;
  rom[03444] = 16'hffff;
  rom[03445] = 16'hffff;
  rom[03446] = 16'hffff;
  rom[03447] = 16'hffff;
  rom[03448] = 16'hffff;
  rom[03449] = 16'hffff;
  rom[03450] = 16'hffff;
  rom[03451] = 16'hffff;
  rom[03452] = 16'hffff;
  rom[03453] = 16'hc618;
  rom[03454] = 16'h3185;
  rom[03455] = 16'h1082;
  rom[03456] = 16'h18c3;
  rom[03457] = 16'h1082;
  rom[03458] = 16'h18c3;
  rom[03459] = 16'h10a2;
  rom[03460] = 16'h18c3;
  rom[03461] = 16'h10a2;
  rom[03462] = 16'h10a2;
  rom[03463] = 16'h10a2;
  rom[03464] = 16'h18e3;
  rom[03465] = 16'h10a2;
  rom[03466] = 16'h18c3;
  rom[03467] = 16'h10a2;
  rom[03468] = 16'h2144;
  rom[03469] = 16'hb616;
  rom[03470] = 16'hfffe;
  rom[03471] = 16'hffff;
  rom[03472] = 16'hffff;
  rom[03473] = 16'hffdf;
  rom[03474] = 16'hffde;
  rom[03475] = 16'h9c8d;
  rom[03476] = 16'hbd4d;
  rom[03477] = 16'hbd0d;
  rom[03478] = 16'h7287;
  rom[03479] = 16'hff7b;
  rom[03480] = 16'hb4af;
  rom[03481] = 16'h7283;
  rom[03482] = 16'hed8e;
  rom[03483] = 16'hf52a;
  rom[03484] = 16'hfd89;
  rom[03485] = 16'hfd48;
  rom[03486] = 16'hf549;
  rom[03487] = 16'hf589;
  rom[03488] = 16'hfe0b;
  rom[03489] = 16'hfd48;
  rom[03490] = 16'hf527;
  rom[03491] = 16'hf568;
  rom[03492] = 16'hfd89;
  rom[03493] = 16'hfd68;
  rom[03494] = 16'hfda9;
  rom[03495] = 16'hfd68;
  rom[03496] = 16'hfd89;
  rom[03497] = 16'hfd68;
  rom[03498] = 16'hfd89;
  rom[03499] = 16'hfd68;
  rom[03500] = 16'hfd89;
  rom[03501] = 16'hfd68;
  rom[03502] = 16'hfd89;
  rom[03503] = 16'hfd88;
  rom[03504] = 16'hfd87;
  rom[03505] = 16'hfd67;
  rom[03506] = 16'hfd69;
  rom[03507] = 16'hfd48;
  rom[03508] = 16'hfd68;
  rom[03509] = 16'hfd67;
  rom[03510] = 16'hfd88;
  rom[03511] = 16'hfd68;
  rom[03512] = 16'hf569;
  rom[03513] = 16'hf569;
  rom[03514] = 16'hf54a;
  rom[03515] = 16'hfdab;
  rom[03516] = 16'he507;
  rom[03517] = 16'hfdc9;
  rom[03518] = 16'hfd47;
  rom[03519] = 16'hfd68;
  rom[03520] = 16'hfd88;
  rom[03521] = 16'hf548;
  rom[03522] = 16'hfdcc;
  rom[03523] = 16'hdd0c;
  rom[03524] = 16'hb44a;
  rom[03525] = 16'h3901;
  rom[03526] = 16'h20c1;
  rom[03527] = 16'h1082;
  rom[03528] = 16'h18a3;
  rom[03529] = 16'h18c3;
  rom[03530] = 16'h18a2;
  rom[03531] = 16'h10a3;
  rom[03532] = 16'h10a3;
  rom[03533] = 16'h10a3;
  rom[03534] = 16'h18a3;
  rom[03535] = 16'h18c3;
  rom[03536] = 16'h1082;
  rom[03537] = 16'h18e3;
  rom[03538] = 16'h1082;
  rom[03539] = 16'h10a2;
  rom[03540] = 16'h7bae;
  rom[03541] = 16'hf77e;
  rom[03542] = 16'hffff;
  rom[03543] = 16'hffff;
  rom[03544] = 16'hffff;
  rom[03545] = 16'hffff;
  rom[03546] = 16'hffff;
  rom[03547] = 16'hffff;
  rom[03548] = 16'hffff;
  rom[03549] = 16'hffff;
  rom[03550] = 16'hffff;
  rom[03551] = 16'hffff;
  rom[03552] = 16'hffff;
  rom[03553] = 16'hffff;
  rom[03554] = 16'hffff;
  rom[03555] = 16'hffff;
  rom[03556] = 16'hffff;
  rom[03557] = 16'hffff;
  rom[03558] = 16'hffff;
  rom[03559] = 16'hffff;
  rom[03560] = 16'hffff;
  rom[03561] = 16'hffff;
  rom[03562] = 16'hffff;
  rom[03563] = 16'hffff;
  rom[03564] = 16'hffff;
  rom[03565] = 16'hffff;
  rom[03566] = 16'hffff;
  rom[03567] = 16'hffff;
  rom[03568] = 16'hffff;
  rom[03569] = 16'hffff;
  rom[03570] = 16'hffff;
  rom[03571] = 16'hffff;
  rom[03572] = 16'hffff;
  rom[03573] = 16'hffff;
  rom[03574] = 16'hffff;
  rom[03575] = 16'hffff;
  rom[03576] = 16'hffff;
  rom[03577] = 16'hffff;
  rom[03578] = 16'hffff;
  rom[03579] = 16'hffff;
  rom[03580] = 16'hffff;
  rom[03581] = 16'hffff;
  rom[03582] = 16'hffff;
  rom[03583] = 16'hffff;
  rom[03584] = 16'hffff;
  rom[03585] = 16'hffff;
  rom[03586] = 16'hffff;
  rom[03587] = 16'hffff;
  rom[03588] = 16'hffff;
  rom[03589] = 16'hffff;
  rom[03590] = 16'hffff;
  rom[03591] = 16'hffff;
  rom[03592] = 16'hffff;
  rom[03593] = 16'hffff;
  rom[03594] = 16'hffff;
  rom[03595] = 16'hffff;
  rom[03596] = 16'hffff;
  rom[03597] = 16'hffff;
  rom[03598] = 16'hffff;
  rom[03599] = 16'hffff;
  rom[03600] = 16'hffff;
  rom[03601] = 16'hffff;
  rom[03602] = 16'hffff;
  rom[03603] = 16'hffff;
  rom[03604] = 16'hffff;
  rom[03605] = 16'hffff;
  rom[03606] = 16'hffff;
  rom[03607] = 16'hffff;
  rom[03608] = 16'hffff;
  rom[03609] = 16'hffff;
  rom[03610] = 16'hffff;
  rom[03611] = 16'hffff;
  rom[03612] = 16'hffff;
  rom[03613] = 16'hffff;
  rom[03614] = 16'hffff;
  rom[03615] = 16'hffff;
  rom[03616] = 16'hffff;
  rom[03617] = 16'hffff;
  rom[03618] = 16'hffff;
  rom[03619] = 16'hffff;
  rom[03620] = 16'hffff;
  rom[03621] = 16'hffff;
  rom[03622] = 16'hffff;
  rom[03623] = 16'hffff;
  rom[03624] = 16'hffff;
  rom[03625] = 16'hffff;
  rom[03626] = 16'hffff;
  rom[03627] = 16'hffff;
  rom[03628] = 16'hffff;
  rom[03629] = 16'hffff;
  rom[03630] = 16'hffff;
  rom[03631] = 16'hffff;
  rom[03632] = 16'hffff;
  rom[03633] = 16'hffff;
  rom[03634] = 16'hffff;
  rom[03635] = 16'hffff;
  rom[03636] = 16'hffff;
  rom[03637] = 16'hffff;
  rom[03638] = 16'hffff;
  rom[03639] = 16'hffff;
  rom[03640] = 16'hffff;
  rom[03641] = 16'hffff;
  rom[03642] = 16'hffff;
  rom[03643] = 16'hffff;
  rom[03644] = 16'hffff;
  rom[03645] = 16'hffff;
  rom[03646] = 16'hffff;
  rom[03647] = 16'hffff;
  rom[03648] = 16'hffff;
  rom[03649] = 16'hffff;
  rom[03650] = 16'hffff;
  rom[03651] = 16'hffff;
  rom[03652] = 16'hffdf;
  rom[03653] = 16'hce39;
  rom[03654] = 16'h2965;
  rom[03655] = 16'h18c3;
  rom[03656] = 16'h1082;
  rom[03657] = 16'h10a2;
  rom[03658] = 16'h18c3;
  rom[03659] = 16'h10a2;
  rom[03660] = 16'h10a2;
  rom[03661] = 16'h10a2;
  rom[03662] = 16'h10a2;
  rom[03663] = 16'h18a3;
  rom[03664] = 16'h18a3;
  rom[03665] = 16'h10a2;
  rom[03666] = 16'h10c2;
  rom[03667] = 16'h18c3;
  rom[03668] = 16'h5b0b;
  rom[03669] = 16'hc658;
  rom[03670] = 16'hef7c;
  rom[03671] = 16'hffdf;
  rom[03672] = 16'hffdf;
  rom[03673] = 16'hffdf;
  rom[03674] = 16'hffbd;
  rom[03675] = 16'h940b;
  rom[03676] = 16'hc52c;
  rom[03677] = 16'hddae;
  rom[03678] = 16'h6203;
  rom[03679] = 16'hb48d;
  rom[03680] = 16'h8326;
  rom[03681] = 16'hc4a9;
  rom[03682] = 16'hedac;
  rom[03683] = 16'hf529;
  rom[03684] = 16'hfd6a;
  rom[03685] = 16'hfd49;
  rom[03686] = 16'hfd68;
  rom[03687] = 16'hfda8;
  rom[03688] = 16'hf546;
  rom[03689] = 16'hfd88;
  rom[03690] = 16'hfd67;
  rom[03691] = 16'hfd89;
  rom[03692] = 16'hfd88;
  rom[03693] = 16'hfd88;
  rom[03694] = 16'hfd68;
  rom[03695] = 16'hfd68;
  rom[03696] = 16'hfd68;
  rom[03697] = 16'hfd88;
  rom[03698] = 16'hf568;
  rom[03699] = 16'hfd88;
  rom[03700] = 16'hfd68;
  rom[03701] = 16'hfd88;
  rom[03702] = 16'hf588;
  rom[03703] = 16'hf5a8;
  rom[03704] = 16'hf587;
  rom[03705] = 16'hfd88;
  rom[03706] = 16'hfd48;
  rom[03707] = 16'hfd68;
  rom[03708] = 16'hfd48;
  rom[03709] = 16'hfd88;
  rom[03710] = 16'hf547;
  rom[03711] = 16'hfd68;
  rom[03712] = 16'hfd68;
  rom[03713] = 16'hfd48;
  rom[03714] = 16'hfd48;
  rom[03715] = 16'hfd69;
  rom[03716] = 16'hf567;
  rom[03717] = 16'hfda8;
  rom[03718] = 16'hf547;
  rom[03719] = 16'hfd88;
  rom[03720] = 16'hf547;
  rom[03721] = 16'hf568;
  rom[03722] = 16'hed49;
  rom[03723] = 16'hed6b;
  rom[03724] = 16'hdd6d;
  rom[03725] = 16'h6a23;
  rom[03726] = 16'h20a0;
  rom[03727] = 16'h18a2;
  rom[03728] = 16'h10a2;
  rom[03729] = 16'h18a3;
  rom[03730] = 16'h18a2;
  rom[03731] = 16'h10a3;
  rom[03732] = 16'h10a3;
  rom[03733] = 16'h10a4;
  rom[03734] = 16'h18a3;
  rom[03735] = 16'h18a3;
  rom[03736] = 16'h18c2;
  rom[03737] = 16'h18c2;
  rom[03738] = 16'h10a1;
  rom[03739] = 16'h18c2;
  rom[03740] = 16'h5aeb;
  rom[03741] = 16'hef3d;
  rom[03742] = 16'hffff;
  rom[03743] = 16'hffff;
  rom[03744] = 16'hffff;
  rom[03745] = 16'hffff;
  rom[03746] = 16'hffff;
  rom[03747] = 16'hffff;
  rom[03748] = 16'hffff;
  rom[03749] = 16'hffff;
  rom[03750] = 16'hffff;
  rom[03751] = 16'hffff;
  rom[03752] = 16'hffff;
  rom[03753] = 16'hffff;
  rom[03754] = 16'hffff;
  rom[03755] = 16'hffff;
  rom[03756] = 16'hffff;
  rom[03757] = 16'hffff;
  rom[03758] = 16'hffff;
  rom[03759] = 16'hffff;
  rom[03760] = 16'hffff;
  rom[03761] = 16'hffff;
  rom[03762] = 16'hffff;
  rom[03763] = 16'hffff;
  rom[03764] = 16'hffff;
  rom[03765] = 16'hffff;
  rom[03766] = 16'hffff;
  rom[03767] = 16'hffff;
  rom[03768] = 16'hffff;
  rom[03769] = 16'hffff;
  rom[03770] = 16'hffff;
  rom[03771] = 16'hffff;
  rom[03772] = 16'hffff;
  rom[03773] = 16'hffff;
  rom[03774] = 16'hffff;
  rom[03775] = 16'hffff;
  rom[03776] = 16'hffff;
  rom[03777] = 16'hffff;
  rom[03778] = 16'hffff;
  rom[03779] = 16'hffff;
  rom[03780] = 16'hffff;
  rom[03781] = 16'hffff;
  rom[03782] = 16'hffff;
  rom[03783] = 16'hffff;
  rom[03784] = 16'hffff;
  rom[03785] = 16'hffff;
  rom[03786] = 16'hffff;
  rom[03787] = 16'hffff;
  rom[03788] = 16'hffff;
  rom[03789] = 16'hffff;
  rom[03790] = 16'hffff;
  rom[03791] = 16'hffff;
  rom[03792] = 16'hffff;
  rom[03793] = 16'hffff;
  rom[03794] = 16'hffff;
  rom[03795] = 16'hffff;
  rom[03796] = 16'hffff;
  rom[03797] = 16'hffff;
  rom[03798] = 16'hffff;
  rom[03799] = 16'hffff;
  rom[03800] = 16'hffff;
  rom[03801] = 16'hffff;
  rom[03802] = 16'hffff;
  rom[03803] = 16'hffff;
  rom[03804] = 16'hffff;
  rom[03805] = 16'hffff;
  rom[03806] = 16'hffff;
  rom[03807] = 16'hffff;
  rom[03808] = 16'hffff;
  rom[03809] = 16'hffff;
  rom[03810] = 16'hffff;
  rom[03811] = 16'hffff;
  rom[03812] = 16'hffff;
  rom[03813] = 16'hffff;
  rom[03814] = 16'hffff;
  rom[03815] = 16'hffff;
  rom[03816] = 16'hffff;
  rom[03817] = 16'hffff;
  rom[03818] = 16'hffff;
  rom[03819] = 16'hffff;
  rom[03820] = 16'hffff;
  rom[03821] = 16'hffff;
  rom[03822] = 16'hffff;
  rom[03823] = 16'hffff;
  rom[03824] = 16'hffff;
  rom[03825] = 16'hffff;
  rom[03826] = 16'hffff;
  rom[03827] = 16'hffff;
  rom[03828] = 16'hffff;
  rom[03829] = 16'hffff;
  rom[03830] = 16'hffff;
  rom[03831] = 16'hffff;
  rom[03832] = 16'hffff;
  rom[03833] = 16'hffff;
  rom[03834] = 16'hffff;
  rom[03835] = 16'hffff;
  rom[03836] = 16'hffff;
  rom[03837] = 16'hffff;
  rom[03838] = 16'hffff;
  rom[03839] = 16'hffff;
  rom[03840] = 16'hffff;
  rom[03841] = 16'hffff;
  rom[03842] = 16'hffff;
  rom[03843] = 16'hffff;
  rom[03844] = 16'hffff;
  rom[03845] = 16'hffff;
  rom[03846] = 16'hffff;
  rom[03847] = 16'hffff;
  rom[03848] = 16'hffff;
  rom[03849] = 16'hffff;
  rom[03850] = 16'hffff;
  rom[03851] = 16'hffff;
  rom[03852] = 16'hffff;
  rom[03853] = 16'hc618;
  rom[03854] = 16'h2965;
  rom[03855] = 16'h18e3;
  rom[03856] = 16'h18a3;
  rom[03857] = 16'h10a2;
  rom[03858] = 16'h18c3;
  rom[03859] = 16'h10a2;
  rom[03860] = 16'h18c3;
  rom[03861] = 16'h10a2;
  rom[03862] = 16'h10a2;
  rom[03863] = 16'h10a2;
  rom[03864] = 16'h18c3;
  rom[03865] = 16'h18c3;
  rom[03866] = 16'h18e3;
  rom[03867] = 16'h18a3;
  rom[03868] = 16'h94b2;
  rom[03869] = 16'h8450;
  rom[03870] = 16'ha534;
  rom[03871] = 16'hff9f;
  rom[03872] = 16'hffff;
  rom[03873] = 16'hff9f;
  rom[03874] = 16'hffbf;
  rom[03875] = 16'h9beb;
  rom[03876] = 16'hd52c;
  rom[03877] = 16'he52c;
  rom[03878] = 16'h9b45;
  rom[03879] = 16'h6a22;
  rom[03880] = 16'hdd4b;
  rom[03881] = 16'hedab;
  rom[03882] = 16'hf56a;
  rom[03883] = 16'hfd6a;
  rom[03884] = 16'hfd6a;
  rom[03885] = 16'hfd69;
  rom[03886] = 16'hfda8;
  rom[03887] = 16'hfd66;
  rom[03888] = 16'hfdc8;
  rom[03889] = 16'hfd88;
  rom[03890] = 16'hfd69;
  rom[03891] = 16'hfd68;
  rom[03892] = 16'hfd69;
  rom[03893] = 16'hfd48;
  rom[03894] = 16'hfd89;
  rom[03895] = 16'hfd68;
  rom[03896] = 16'hfd89;
  rom[03897] = 16'hfd68;
  rom[03898] = 16'hfd89;
  rom[03899] = 16'hfd68;
  rom[03900] = 16'hfd89;
  rom[03901] = 16'hfd88;
  rom[03902] = 16'hfda9;
  rom[03903] = 16'hf588;
  rom[03904] = 16'hf5a9;
  rom[03905] = 16'hfd88;
  rom[03906] = 16'hfd89;
  rom[03907] = 16'hfd48;
  rom[03908] = 16'hfd69;
  rom[03909] = 16'hfd68;
  rom[03910] = 16'hfd87;
  rom[03911] = 16'hfd47;
  rom[03912] = 16'hfd89;
  rom[03913] = 16'hfd48;
  rom[03914] = 16'hfd89;
  rom[03915] = 16'hfd47;
  rom[03916] = 16'hfd67;
  rom[03917] = 16'hfd88;
  rom[03918] = 16'hfd89;
  rom[03919] = 16'hf548;
  rom[03920] = 16'hfd89;
  rom[03921] = 16'hf567;
  rom[03922] = 16'hfda9;
  rom[03923] = 16'hf529;
  rom[03924] = 16'he56c;
  rom[03925] = 16'ha3e9;
  rom[03926] = 16'h3902;
  rom[03927] = 16'h1881;
  rom[03928] = 16'h18e3;
  rom[03929] = 16'h10a2;
  rom[03930] = 16'h18a2;
  rom[03931] = 16'h10a3;
  rom[03932] = 16'h10a4;
  rom[03933] = 16'h10a4;
  rom[03934] = 16'h18a3;
  rom[03935] = 16'h18a2;
  rom[03936] = 16'h18c2;
  rom[03937] = 16'h1082;
  rom[03938] = 16'h2103;
  rom[03939] = 16'h10a2;
  rom[03940] = 16'h5acb;
  rom[03941] = 16'hef3d;
  rom[03942] = 16'hffff;
  rom[03943] = 16'hffff;
  rom[03944] = 16'hffff;
  rom[03945] = 16'hffff;
  rom[03946] = 16'hffff;
  rom[03947] = 16'hffff;
  rom[03948] = 16'hffff;
  rom[03949] = 16'hffff;
  rom[03950] = 16'hffff;
  rom[03951] = 16'hffff;
  rom[03952] = 16'hffff;
  rom[03953] = 16'hffff;
  rom[03954] = 16'hffff;
  rom[03955] = 16'hffff;
  rom[03956] = 16'hffff;
  rom[03957] = 16'hffff;
  rom[03958] = 16'hffff;
  rom[03959] = 16'hffff;
  rom[03960] = 16'hffff;
  rom[03961] = 16'hffff;
  rom[03962] = 16'hffff;
  rom[03963] = 16'hffff;
  rom[03964] = 16'hffff;
  rom[03965] = 16'hffff;
  rom[03966] = 16'hffff;
  rom[03967] = 16'hffff;
  rom[03968] = 16'hffff;
  rom[03969] = 16'hffff;
  rom[03970] = 16'hffff;
  rom[03971] = 16'hffff;
  rom[03972] = 16'hffff;
  rom[03973] = 16'hffff;
  rom[03974] = 16'hffff;
  rom[03975] = 16'hffff;
  rom[03976] = 16'hffff;
  rom[03977] = 16'hffff;
  rom[03978] = 16'hffff;
  rom[03979] = 16'hffff;
  rom[03980] = 16'hffff;
  rom[03981] = 16'hffff;
  rom[03982] = 16'hffff;
  rom[03983] = 16'hffff;
  rom[03984] = 16'hffff;
  rom[03985] = 16'hffff;
  rom[03986] = 16'hffff;
  rom[03987] = 16'hffff;
  rom[03988] = 16'hffff;
  rom[03989] = 16'hffff;
  rom[03990] = 16'hffff;
  rom[03991] = 16'hffff;
  rom[03992] = 16'hffff;
  rom[03993] = 16'hffff;
  rom[03994] = 16'hffff;
  rom[03995] = 16'hffff;
  rom[03996] = 16'hffff;
  rom[03997] = 16'hffff;
  rom[03998] = 16'hffff;
  rom[03999] = 16'hffff;
  rom[04000] = 16'hffff;
  rom[04001] = 16'hffff;
  rom[04002] = 16'hffff;
  rom[04003] = 16'hffff;
  rom[04004] = 16'hffff;
  rom[04005] = 16'hffff;
  rom[04006] = 16'hffff;
  rom[04007] = 16'hffff;
  rom[04008] = 16'hffff;
  rom[04009] = 16'hffff;
  rom[04010] = 16'hffff;
  rom[04011] = 16'hffff;
  rom[04012] = 16'hffff;
  rom[04013] = 16'hffff;
  rom[04014] = 16'hffff;
  rom[04015] = 16'hffff;
  rom[04016] = 16'hffff;
  rom[04017] = 16'hffff;
  rom[04018] = 16'hffff;
  rom[04019] = 16'hffff;
  rom[04020] = 16'hffff;
  rom[04021] = 16'hffff;
  rom[04022] = 16'hffff;
  rom[04023] = 16'hffff;
  rom[04024] = 16'hffff;
  rom[04025] = 16'hffff;
  rom[04026] = 16'hffff;
  rom[04027] = 16'hffff;
  rom[04028] = 16'hffff;
  rom[04029] = 16'hffff;
  rom[04030] = 16'hffff;
  rom[04031] = 16'hffff;
  rom[04032] = 16'hffff;
  rom[04033] = 16'hffff;
  rom[04034] = 16'hffff;
  rom[04035] = 16'hffff;
  rom[04036] = 16'hffff;
  rom[04037] = 16'hffff;
  rom[04038] = 16'hffff;
  rom[04039] = 16'hffff;
  rom[04040] = 16'hffff;
  rom[04041] = 16'hffff;
  rom[04042] = 16'hffff;
  rom[04043] = 16'hffff;
  rom[04044] = 16'hffff;
  rom[04045] = 16'hffff;
  rom[04046] = 16'hffff;
  rom[04047] = 16'hffff;
  rom[04048] = 16'hffff;
  rom[04049] = 16'hffff;
  rom[04050] = 16'hffff;
  rom[04051] = 16'hffff;
  rom[04052] = 16'hffff;
  rom[04053] = 16'hc618;
  rom[04054] = 16'h2965;
  rom[04055] = 16'h10a2;
  rom[04056] = 16'h10a2;
  rom[04057] = 16'h10a2;
  rom[04058] = 16'h10a2;
  rom[04059] = 16'h10a2;
  rom[04060] = 16'h10a2;
  rom[04061] = 16'h10a2;
  rom[04062] = 16'h10a2;
  rom[04063] = 16'h10a2;
  rom[04064] = 16'h10a2;
  rom[04065] = 16'h18c3;
  rom[04066] = 16'h10c2;
  rom[04067] = 16'h3166;
  rom[04068] = 16'hbdf7;
  rom[04069] = 16'hc637;
  rom[04070] = 16'h5b0b;
  rom[04071] = 16'hde7a;
  rom[04072] = 16'hff7e;
  rom[04073] = 16'hffbf;
  rom[04074] = 16'hde57;
  rom[04075] = 16'h8b27;
  rom[04076] = 16'hdd4b;
  rom[04077] = 16'hf58b;
  rom[04078] = 16'he50a;
  rom[04079] = 16'hd4e9;
  rom[04080] = 16'he5aa;
  rom[04081] = 16'hed89;
  rom[04082] = 16'hf568;
  rom[04083] = 16'hfda9;
  rom[04084] = 16'hf548;
  rom[04085] = 16'hfd89;
  rom[04086] = 16'hf587;
  rom[04087] = 16'hfda8;
  rom[04088] = 16'hf587;
  rom[04089] = 16'hfd89;
  rom[04090] = 16'hfd68;
  rom[04091] = 16'hfd89;
  rom[04092] = 16'hf568;
  rom[04093] = 16'hfd89;
  rom[04094] = 16'hfd88;
  rom[04095] = 16'hfd88;
  rom[04096] = 16'hf588;
  rom[04097] = 16'hfd88;
  rom[04098] = 16'hfd68;
  rom[04099] = 16'hfd88;
  rom[04100] = 16'hf568;
  rom[04101] = 16'hfd88;
  rom[04102] = 16'hfd88;
  rom[04103] = 16'hf5a8;
  rom[04104] = 16'hf588;
  rom[04105] = 16'hfda8;
  rom[04106] = 16'hfd68;
  rom[04107] = 16'hfd88;
  rom[04108] = 16'hf568;
  rom[04109] = 16'hfd88;
  rom[04110] = 16'hfd68;
  rom[04111] = 16'hfd68;
  rom[04112] = 16'hfd47;
  rom[04113] = 16'hfd68;
  rom[04114] = 16'hfd48;
  rom[04115] = 16'hfd68;
  rom[04116] = 16'hfd88;
  rom[04117] = 16'hf548;
  rom[04118] = 16'hf549;
  rom[04119] = 16'hfdaa;
  rom[04120] = 16'hf567;
  rom[04121] = 16'hfd87;
  rom[04122] = 16'hf567;
  rom[04123] = 16'hfd49;
  rom[04124] = 16'hed6b;
  rom[04125] = 16'hb44a;
  rom[04126] = 16'h3101;
  rom[04127] = 16'h18a2;
  rom[04128] = 16'h1082;
  rom[04129] = 16'h18c2;
  rom[04130] = 16'h18a2;
  rom[04131] = 16'h10a2;
  rom[04132] = 16'h10a3;
  rom[04133] = 16'h10a3;
  rom[04134] = 16'h18a2;
  rom[04135] = 16'h18c2;
  rom[04136] = 16'h1082;
  rom[04137] = 16'h18a2;
  rom[04138] = 16'h18c2;
  rom[04139] = 16'h10a2;
  rom[04140] = 16'h632c;
  rom[04141] = 16'hf77e;
  rom[04142] = 16'hffff;
  rom[04143] = 16'hffff;
  rom[04144] = 16'hffff;
  rom[04145] = 16'hffff;
  rom[04146] = 16'hffff;
  rom[04147] = 16'hffff;
  rom[04148] = 16'hffff;
  rom[04149] = 16'hffff;
  rom[04150] = 16'hffff;
  rom[04151] = 16'hffff;
  rom[04152] = 16'hffff;
  rom[04153] = 16'hffff;
  rom[04154] = 16'hffff;
  rom[04155] = 16'hffff;
  rom[04156] = 16'hffff;
  rom[04157] = 16'hffff;
  rom[04158] = 16'hffff;
  rom[04159] = 16'hffff;
  rom[04160] = 16'hffff;
  rom[04161] = 16'hffff;
  rom[04162] = 16'hffff;
  rom[04163] = 16'hffff;
  rom[04164] = 16'hffff;
  rom[04165] = 16'hffff;
  rom[04166] = 16'hffff;
  rom[04167] = 16'hffff;
  rom[04168] = 16'hffff;
  rom[04169] = 16'hffff;
  rom[04170] = 16'hffff;
  rom[04171] = 16'hffff;
  rom[04172] = 16'hffff;
  rom[04173] = 16'hffff;
  rom[04174] = 16'hffff;
  rom[04175] = 16'hffff;
  rom[04176] = 16'hffff;
  rom[04177] = 16'hffff;
  rom[04178] = 16'hffff;
  rom[04179] = 16'hffff;
  rom[04180] = 16'hffff;
  rom[04181] = 16'hffff;
  rom[04182] = 16'hffff;
  rom[04183] = 16'hffff;
  rom[04184] = 16'hffff;
  rom[04185] = 16'hffff;
  rom[04186] = 16'hffff;
  rom[04187] = 16'hffff;
  rom[04188] = 16'hffff;
  rom[04189] = 16'hffff;
  rom[04190] = 16'hffff;
  rom[04191] = 16'hffff;
  rom[04192] = 16'hffff;
  rom[04193] = 16'hffff;
  rom[04194] = 16'hffff;
  rom[04195] = 16'hffff;
  rom[04196] = 16'hffff;
  rom[04197] = 16'hffff;
  rom[04198] = 16'hffff;
  rom[04199] = 16'hffff;
  rom[04200] = 16'hffff;
  rom[04201] = 16'hffff;
  rom[04202] = 16'hffff;
  rom[04203] = 16'hffff;
  rom[04204] = 16'hffff;
  rom[04205] = 16'hffff;
  rom[04206] = 16'hffff;
  rom[04207] = 16'hffff;
  rom[04208] = 16'hffff;
  rom[04209] = 16'hffff;
  rom[04210] = 16'hffff;
  rom[04211] = 16'hffff;
  rom[04212] = 16'hffff;
  rom[04213] = 16'hffff;
  rom[04214] = 16'hffff;
  rom[04215] = 16'hffff;
  rom[04216] = 16'hffff;
  rom[04217] = 16'hffff;
  rom[04218] = 16'hffff;
  rom[04219] = 16'hffff;
  rom[04220] = 16'hffff;
  rom[04221] = 16'hffff;
  rom[04222] = 16'hffff;
  rom[04223] = 16'hffff;
  rom[04224] = 16'hffff;
  rom[04225] = 16'hffff;
  rom[04226] = 16'hffff;
  rom[04227] = 16'hffff;
  rom[04228] = 16'hffff;
  rom[04229] = 16'hffff;
  rom[04230] = 16'hffff;
  rom[04231] = 16'hffff;
  rom[04232] = 16'hffff;
  rom[04233] = 16'hffff;
  rom[04234] = 16'hffff;
  rom[04235] = 16'hffff;
  rom[04236] = 16'hffff;
  rom[04237] = 16'hffff;
  rom[04238] = 16'hffff;
  rom[04239] = 16'hffff;
  rom[04240] = 16'hffff;
  rom[04241] = 16'hffff;
  rom[04242] = 16'hffff;
  rom[04243] = 16'hffff;
  rom[04244] = 16'hffff;
  rom[04245] = 16'hffff;
  rom[04246] = 16'hffff;
  rom[04247] = 16'hffff;
  rom[04248] = 16'hffff;
  rom[04249] = 16'hffff;
  rom[04250] = 16'hffff;
  rom[04251] = 16'hffff;
  rom[04252] = 16'hffff;
  rom[04253] = 16'hc618;
  rom[04254] = 16'h3185;
  rom[04255] = 16'h10a2;
  rom[04256] = 16'h18e3;
  rom[04257] = 16'h10a2;
  rom[04258] = 16'h18c3;
  rom[04259] = 16'h10a2;
  rom[04260] = 16'h18c3;
  rom[04261] = 16'h10a2;
  rom[04262] = 16'h18c3;
  rom[04263] = 16'h10a2;
  rom[04264] = 16'h1082;
  rom[04265] = 16'h18c3;
  rom[04266] = 16'h18a3;
  rom[04267] = 16'h4a28;
  rom[04268] = 16'he6fc;
  rom[04269] = 16'hef5c;
  rom[04270] = 16'h6b0b;
  rom[04271] = 16'h6aeb;
  rom[04272] = 16'he699;
  rom[04273] = 16'hff7c;
  rom[04274] = 16'hb4b0;
  rom[04275] = 16'habc9;
  rom[04276] = 16'hed4a;
  rom[04277] = 16'hfda9;
  rom[04278] = 16'hf569;
  rom[04279] = 16'hedaa;
  rom[04280] = 16'hf5ca;
  rom[04281] = 16'hed67;
  rom[04282] = 16'hfda8;
  rom[04283] = 16'hf587;
  rom[04284] = 16'hfda9;
  rom[04285] = 16'hf5a9;
  rom[04286] = 16'hf5a9;
  rom[04287] = 16'hf588;
  rom[04288] = 16'hfda9;
  rom[04289] = 16'hfd69;
  rom[04290] = 16'hfdaa;
  rom[04291] = 16'hfd8a;
  rom[04292] = 16'hfd89;
  rom[04293] = 16'hfd88;
  rom[04294] = 16'hfd89;
  rom[04295] = 16'hfd88;
  rom[04296] = 16'hfda9;
  rom[04297] = 16'hfd88;
  rom[04298] = 16'hfda9;
  rom[04299] = 16'hfd88;
  rom[04300] = 16'hfda9;
  rom[04301] = 16'hfd69;
  rom[04302] = 16'hfd8a;
  rom[04303] = 16'hfd89;
  rom[04304] = 16'hfda9;
  rom[04305] = 16'hfd88;
  rom[04306] = 16'hfd89;
  rom[04307] = 16'hfd88;
  rom[04308] = 16'hfda9;
  rom[04309] = 16'hf588;
  rom[04310] = 16'hfd89;
  rom[04311] = 16'hfd68;
  rom[04312] = 16'hfd68;
  rom[04313] = 16'hfd88;
  rom[04314] = 16'hfd69;
  rom[04315] = 16'hfd89;
  rom[04316] = 16'hfd69;
  rom[04317] = 16'hfd4a;
  rom[04318] = 16'hfd6b;
  rom[04319] = 16'hfd69;
  rom[04320] = 16'hfd88;
  rom[04321] = 16'hfd86;
  rom[04322] = 16'hfd67;
  rom[04323] = 16'hfd68;
  rom[04324] = 16'hed4a;
  rom[04325] = 16'hcceb;
  rom[04326] = 16'h51a4;
  rom[04327] = 16'h20a2;
  rom[04328] = 16'h18a3;
  rom[04329] = 16'h18c2;
  rom[04330] = 16'h18c2;
  rom[04331] = 16'h10a2;
  rom[04332] = 16'h10a3;
  rom[04333] = 16'h10a3;
  rom[04334] = 16'h18a3;
  rom[04335] = 16'h18a2;
  rom[04336] = 16'h18a2;
  rom[04337] = 16'h10a2;
  rom[04338] = 16'h18c2;
  rom[04339] = 16'h10a2;
  rom[04340] = 16'h7bae;
  rom[04341] = 16'hf79e;
  rom[04342] = 16'hffff;
  rom[04343] = 16'hffff;
  rom[04344] = 16'hffff;
  rom[04345] = 16'hffff;
  rom[04346] = 16'hffff;
  rom[04347] = 16'hffff;
  rom[04348] = 16'hffff;
  rom[04349] = 16'hffff;
  rom[04350] = 16'hffff;
  rom[04351] = 16'hffff;
  rom[04352] = 16'hffff;
  rom[04353] = 16'hffff;
  rom[04354] = 16'hffff;
  rom[04355] = 16'hffff;
  rom[04356] = 16'hffff;
  rom[04357] = 16'hffff;
  rom[04358] = 16'hffff;
  rom[04359] = 16'hffff;
  rom[04360] = 16'hffff;
  rom[04361] = 16'hffff;
  rom[04362] = 16'hffff;
  rom[04363] = 16'hffff;
  rom[04364] = 16'hffff;
  rom[04365] = 16'hffff;
  rom[04366] = 16'hffff;
  rom[04367] = 16'hffff;
  rom[04368] = 16'hffff;
  rom[04369] = 16'hffff;
  rom[04370] = 16'hffff;
  rom[04371] = 16'hffff;
  rom[04372] = 16'hffff;
  rom[04373] = 16'hffff;
  rom[04374] = 16'hffff;
  rom[04375] = 16'hffff;
  rom[04376] = 16'hffff;
  rom[04377] = 16'hffff;
  rom[04378] = 16'hffff;
  rom[04379] = 16'hffff;
  rom[04380] = 16'hffff;
  rom[04381] = 16'hffff;
  rom[04382] = 16'hffff;
  rom[04383] = 16'hffff;
  rom[04384] = 16'hffff;
  rom[04385] = 16'hffff;
  rom[04386] = 16'hffff;
  rom[04387] = 16'hffff;
  rom[04388] = 16'hffff;
  rom[04389] = 16'hffff;
  rom[04390] = 16'hffff;
  rom[04391] = 16'hffff;
  rom[04392] = 16'hffff;
  rom[04393] = 16'hffff;
  rom[04394] = 16'hffff;
  rom[04395] = 16'hffff;
  rom[04396] = 16'hffff;
  rom[04397] = 16'hffff;
  rom[04398] = 16'hffff;
  rom[04399] = 16'hffff;
  rom[04400] = 16'hffff;
  rom[04401] = 16'hffff;
  rom[04402] = 16'hffff;
  rom[04403] = 16'hffff;
  rom[04404] = 16'hffff;
  rom[04405] = 16'hffff;
  rom[04406] = 16'hffff;
  rom[04407] = 16'hffff;
  rom[04408] = 16'hffff;
  rom[04409] = 16'hffff;
  rom[04410] = 16'hffff;
  rom[04411] = 16'hffff;
  rom[04412] = 16'hffff;
  rom[04413] = 16'hffff;
  rom[04414] = 16'hffff;
  rom[04415] = 16'hffff;
  rom[04416] = 16'hffff;
  rom[04417] = 16'hffff;
  rom[04418] = 16'hffff;
  rom[04419] = 16'hffff;
  rom[04420] = 16'hffff;
  rom[04421] = 16'hffff;
  rom[04422] = 16'hffff;
  rom[04423] = 16'hffff;
  rom[04424] = 16'hffff;
  rom[04425] = 16'hffff;
  rom[04426] = 16'hffff;
  rom[04427] = 16'hffff;
  rom[04428] = 16'hffff;
  rom[04429] = 16'hffff;
  rom[04430] = 16'hffff;
  rom[04431] = 16'hffff;
  rom[04432] = 16'hffff;
  rom[04433] = 16'hffff;
  rom[04434] = 16'hffff;
  rom[04435] = 16'hffff;
  rom[04436] = 16'hffff;
  rom[04437] = 16'hffff;
  rom[04438] = 16'hffff;
  rom[04439] = 16'hffff;
  rom[04440] = 16'hffff;
  rom[04441] = 16'hffff;
  rom[04442] = 16'hffff;
  rom[04443] = 16'hffff;
  rom[04444] = 16'hffff;
  rom[04445] = 16'hffff;
  rom[04446] = 16'hffff;
  rom[04447] = 16'hffff;
  rom[04448] = 16'hffff;
  rom[04449] = 16'hffff;
  rom[04450] = 16'hffff;
  rom[04451] = 16'hffff;
  rom[04452] = 16'hffff;
  rom[04453] = 16'hd679;
  rom[04454] = 16'h3185;
  rom[04455] = 16'h18c2;
  rom[04456] = 16'h18c2;
  rom[04457] = 16'h10a2;
  rom[04458] = 16'h10a2;
  rom[04459] = 16'h10a2;
  rom[04460] = 16'h10a3;
  rom[04461] = 16'h18c3;
  rom[04462] = 16'h10a2;
  rom[04463] = 16'h18c3;
  rom[04464] = 16'h0861;
  rom[04465] = 16'h18e3;
  rom[04466] = 16'h0861;
  rom[04467] = 16'h526a;
  rom[04468] = 16'hef3c;
  rom[04469] = 16'hfffe;
  rom[04470] = 16'h840d;
  rom[04471] = 16'h62a8;
  rom[04472] = 16'h8369;
  rom[04473] = 16'hb4ae;
  rom[04474] = 16'h6a02;
  rom[04475] = 16'hd4ea;
  rom[04476] = 16'hed48;
  rom[04477] = 16'hfd88;
  rom[04478] = 16'hfd68;
  rom[04479] = 16'hf5aa;
  rom[04480] = 16'hf588;
  rom[04481] = 16'hfda8;
  rom[04482] = 16'hf587;
  rom[04483] = 16'hfda8;
  rom[04484] = 16'hf587;
  rom[04485] = 16'hf5a8;
  rom[04486] = 16'hf588;
  rom[04487] = 16'hfda9;
  rom[04488] = 16'hf568;
  rom[04489] = 16'hfd8a;
  rom[04490] = 16'hf589;
  rom[04491] = 16'hf589;
  rom[04492] = 16'hfd89;
  rom[04493] = 16'hfda9;
  rom[04494] = 16'hf588;
  rom[04495] = 16'hfda8;
  rom[04496] = 16'hfd88;
  rom[04497] = 16'hfda8;
  rom[04498] = 16'hf588;
  rom[04499] = 16'hfda9;
  rom[04500] = 16'hfd89;
  rom[04501] = 16'hfd89;
  rom[04502] = 16'hfd69;
  rom[04503] = 16'hfd88;
  rom[04504] = 16'hfd88;
  rom[04505] = 16'hfda8;
  rom[04506] = 16'hf588;
  rom[04507] = 16'hfda8;
  rom[04508] = 16'hf588;
  rom[04509] = 16'hf5a8;
  rom[04510] = 16'hf568;
  rom[04511] = 16'hfd88;
  rom[04512] = 16'hfd68;
  rom[04513] = 16'hfda8;
  rom[04514] = 16'hf589;
  rom[04515] = 16'hf549;
  rom[04516] = 16'hfd49;
  rom[04517] = 16'hfd6a;
  rom[04518] = 16'hf549;
  rom[04519] = 16'hfd89;
  rom[04520] = 16'hf547;
  rom[04521] = 16'hfd87;
  rom[04522] = 16'hf566;
  rom[04523] = 16'hfd69;
  rom[04524] = 16'hf56a;
  rom[04525] = 16'hd50d;
  rom[04526] = 16'h5a05;
  rom[04527] = 16'h20a2;
  rom[04528] = 16'h18a2;
  rom[04529] = 16'h18e3;
  rom[04530] = 16'h10a1;
  rom[04531] = 16'h10c2;
  rom[04532] = 16'h10a2;
  rom[04533] = 16'h10a3;
  rom[04534] = 16'h10a2;
  rom[04535] = 16'h18a2;
  rom[04536] = 16'h10a2;
  rom[04537] = 16'h18a2;
  rom[04538] = 16'h10a2;
  rom[04539] = 16'h10a2;
  rom[04540] = 16'h73ae;
  rom[04541] = 16'hffbf;
  rom[04542] = 16'hffff;
  rom[04543] = 16'hffff;
  rom[04544] = 16'hffff;
  rom[04545] = 16'hffff;
  rom[04546] = 16'hffff;
  rom[04547] = 16'hffff;
  rom[04548] = 16'hffff;
  rom[04549] = 16'hffff;
  rom[04550] = 16'hffff;
  rom[04551] = 16'hffff;
  rom[04552] = 16'hffff;
  rom[04553] = 16'hffff;
  rom[04554] = 16'hffff;
  rom[04555] = 16'hffff;
  rom[04556] = 16'hffff;
  rom[04557] = 16'hffff;
  rom[04558] = 16'hffff;
  rom[04559] = 16'hffff;
  rom[04560] = 16'hffff;
  rom[04561] = 16'hffff;
  rom[04562] = 16'hffff;
  rom[04563] = 16'hffff;
  rom[04564] = 16'hffff;
  rom[04565] = 16'hffff;
  rom[04566] = 16'hffff;
  rom[04567] = 16'hffff;
  rom[04568] = 16'hffff;
  rom[04569] = 16'hffff;
  rom[04570] = 16'hffff;
  rom[04571] = 16'hffff;
  rom[04572] = 16'hffff;
  rom[04573] = 16'hffff;
  rom[04574] = 16'hffff;
  rom[04575] = 16'hffff;
  rom[04576] = 16'hffff;
  rom[04577] = 16'hffff;
  rom[04578] = 16'hffff;
  rom[04579] = 16'hffff;
  rom[04580] = 16'hffff;
  rom[04581] = 16'hffff;
  rom[04582] = 16'hffff;
  rom[04583] = 16'hffff;
  rom[04584] = 16'hffff;
  rom[04585] = 16'hffff;
  rom[04586] = 16'hffff;
  rom[04587] = 16'hffff;
  rom[04588] = 16'hffff;
  rom[04589] = 16'hffff;
  rom[04590] = 16'hffff;
  rom[04591] = 16'hffff;
  rom[04592] = 16'hffff;
  rom[04593] = 16'hffff;
  rom[04594] = 16'hffff;
  rom[04595] = 16'hffff;
  rom[04596] = 16'hffff;
  rom[04597] = 16'hffff;
  rom[04598] = 16'hffff;
  rom[04599] = 16'hffff;
  rom[04600] = 16'hffff;
  rom[04601] = 16'hffff;
  rom[04602] = 16'hffff;
  rom[04603] = 16'hffff;
  rom[04604] = 16'hffff;
  rom[04605] = 16'hffff;
  rom[04606] = 16'hffff;
  rom[04607] = 16'hffff;
  rom[04608] = 16'hffff;
  rom[04609] = 16'hffff;
  rom[04610] = 16'hffff;
  rom[04611] = 16'hffff;
  rom[04612] = 16'hffff;
  rom[04613] = 16'hffff;
  rom[04614] = 16'hffff;
  rom[04615] = 16'hffff;
  rom[04616] = 16'hffff;
  rom[04617] = 16'hffff;
  rom[04618] = 16'hffff;
  rom[04619] = 16'hffff;
  rom[04620] = 16'hffff;
  rom[04621] = 16'hffff;
  rom[04622] = 16'hffff;
  rom[04623] = 16'hffff;
  rom[04624] = 16'hffff;
  rom[04625] = 16'hffff;
  rom[04626] = 16'hffff;
  rom[04627] = 16'hffff;
  rom[04628] = 16'hffff;
  rom[04629] = 16'hffff;
  rom[04630] = 16'hffff;
  rom[04631] = 16'hffff;
  rom[04632] = 16'hffff;
  rom[04633] = 16'hffff;
  rom[04634] = 16'hffff;
  rom[04635] = 16'hffff;
  rom[04636] = 16'hffff;
  rom[04637] = 16'hffff;
  rom[04638] = 16'hffff;
  rom[04639] = 16'hffff;
  rom[04640] = 16'hffff;
  rom[04641] = 16'hffff;
  rom[04642] = 16'hffff;
  rom[04643] = 16'hffff;
  rom[04644] = 16'hffff;
  rom[04645] = 16'hffff;
  rom[04646] = 16'hffff;
  rom[04647] = 16'hffff;
  rom[04648] = 16'hffff;
  rom[04649] = 16'hffff;
  rom[04650] = 16'hffff;
  rom[04651] = 16'hffff;
  rom[04652] = 16'hffff;
  rom[04653] = 16'hd69a;
  rom[04654] = 16'h39c7;
  rom[04655] = 16'h18c2;
  rom[04656] = 16'h18c2;
  rom[04657] = 16'h10c2;
  rom[04658] = 16'h18a3;
  rom[04659] = 16'h18a3;
  rom[04660] = 16'h10a3;
  rom[04661] = 16'h18a3;
  rom[04662] = 16'h10c2;
  rom[04663] = 16'h10c2;
  rom[04664] = 16'h10a2;
  rom[04665] = 16'h10a2;
  rom[04666] = 16'h20c4;
  rom[04667] = 16'h526a;
  rom[04668] = 16'hf77e;
  rom[04669] = 16'hffde;
  rom[04670] = 16'hb512;
  rom[04671] = 16'h9c0c;
  rom[04672] = 16'hc4cd;
  rom[04673] = 16'ha3c8;
  rom[04674] = 16'hccca;
  rom[04675] = 16'he549;
  rom[04676] = 16'hfdc9;
  rom[04677] = 16'hf546;
  rom[04678] = 16'hfd89;
  rom[04679] = 16'hfd89;
  rom[04680] = 16'hfd89;
  rom[04681] = 16'hfd88;
  rom[04682] = 16'hfda9;
  rom[04683] = 16'hfd88;
  rom[04684] = 16'hfd88;
  rom[04685] = 16'hfd88;
  rom[04686] = 16'hfda9;
  rom[04687] = 16'hfd88;
  rom[04688] = 16'hfda9;
  rom[04689] = 16'hfd89;
  rom[04690] = 16'hfda9;
  rom[04691] = 16'hfd88;
  rom[04692] = 16'hfda9;
  rom[04693] = 16'hfd88;
  rom[04694] = 16'hfda9;
  rom[04695] = 16'hfd88;
  rom[04696] = 16'hfda9;
  rom[04697] = 16'hfd88;
  rom[04698] = 16'hfda9;
  rom[04699] = 16'hfd88;
  rom[04700] = 16'hfda9;
  rom[04701] = 16'hfd88;
  rom[04702] = 16'hfda9;
  rom[04703] = 16'hfd88;
  rom[04704] = 16'hfda9;
  rom[04705] = 16'hfd88;
  rom[04706] = 16'hfda9;
  rom[04707] = 16'hfda8;
  rom[04708] = 16'hfda9;
  rom[04709] = 16'hfd88;
  rom[04710] = 16'hfda9;
  rom[04711] = 16'hfd88;
  rom[04712] = 16'hfda9;
  rom[04713] = 16'hf5a8;
  rom[04714] = 16'hfd89;
  rom[04715] = 16'hfd69;
  rom[04716] = 16'hfd6a;
  rom[04717] = 16'hfd89;
  rom[04718] = 16'hfd89;
  rom[04719] = 16'hfd88;
  rom[04720] = 16'hfd68;
  rom[04721] = 16'hfd68;
  rom[04722] = 16'hfd68;
  rom[04723] = 16'hfd69;
  rom[04724] = 16'hfd8a;
  rom[04725] = 16'hd50d;
  rom[04726] = 16'h6206;
  rom[04727] = 16'h1881;
  rom[04728] = 16'h20a3;
  rom[04729] = 16'h18a2;
  rom[04730] = 16'h10c2;
  rom[04731] = 16'h10e2;
  rom[04732] = 16'h10a3;
  rom[04733] = 16'h10a3;
  rom[04734] = 16'h10c3;
  rom[04735] = 16'h10a2;
  rom[04736] = 16'h18c2;
  rom[04737] = 16'h18a2;
  rom[04738] = 16'h10a2;
  rom[04739] = 16'h18a2;
  rom[04740] = 16'h8c11;
  rom[04741] = 16'hffdf;
  rom[04742] = 16'hffff;
  rom[04743] = 16'hffff;
  rom[04744] = 16'hffff;
  rom[04745] = 16'hffff;
  rom[04746] = 16'hffff;
  rom[04747] = 16'hffff;
  rom[04748] = 16'hffff;
  rom[04749] = 16'hffff;
  rom[04750] = 16'hffff;
  rom[04751] = 16'hffff;
  rom[04752] = 16'hffff;
  rom[04753] = 16'hffff;
  rom[04754] = 16'hffff;
  rom[04755] = 16'hffff;
  rom[04756] = 16'hffff;
  rom[04757] = 16'hffff;
  rom[04758] = 16'hffff;
  rom[04759] = 16'hffff;
  rom[04760] = 16'hffff;
  rom[04761] = 16'hffff;
  rom[04762] = 16'hffff;
  rom[04763] = 16'hffff;
  rom[04764] = 16'hffff;
  rom[04765] = 16'hffff;
  rom[04766] = 16'hffff;
  rom[04767] = 16'hffff;
  rom[04768] = 16'hffff;
  rom[04769] = 16'hffff;
  rom[04770] = 16'hffff;
  rom[04771] = 16'hffff;
  rom[04772] = 16'hffff;
  rom[04773] = 16'hffff;
  rom[04774] = 16'hffff;
  rom[04775] = 16'hffff;
  rom[04776] = 16'hffff;
  rom[04777] = 16'hffff;
  rom[04778] = 16'hffff;
  rom[04779] = 16'hffff;
  rom[04780] = 16'hffff;
  rom[04781] = 16'hffff;
  rom[04782] = 16'hffff;
  rom[04783] = 16'hffff;
  rom[04784] = 16'hffff;
  rom[04785] = 16'hffff;
  rom[04786] = 16'hffff;
  rom[04787] = 16'hffff;
  rom[04788] = 16'hffff;
  rom[04789] = 16'hffff;
  rom[04790] = 16'hffff;
  rom[04791] = 16'hffff;
  rom[04792] = 16'hffff;
  rom[04793] = 16'hffff;
  rom[04794] = 16'hffff;
  rom[04795] = 16'hffff;
  rom[04796] = 16'hffff;
  rom[04797] = 16'hffff;
  rom[04798] = 16'hffff;
  rom[04799] = 16'hffff;
  rom[04800] = 16'hffff;
  rom[04801] = 16'hffff;
  rom[04802] = 16'hffff;
  rom[04803] = 16'hffff;
  rom[04804] = 16'hffff;
  rom[04805] = 16'hffff;
  rom[04806] = 16'hffff;
  rom[04807] = 16'hffff;
  rom[04808] = 16'hffff;
  rom[04809] = 16'hffff;
  rom[04810] = 16'hffff;
  rom[04811] = 16'hffff;
  rom[04812] = 16'hffff;
  rom[04813] = 16'hffff;
  rom[04814] = 16'hffff;
  rom[04815] = 16'hffff;
  rom[04816] = 16'hffff;
  rom[04817] = 16'hffff;
  rom[04818] = 16'hffff;
  rom[04819] = 16'hffff;
  rom[04820] = 16'hffff;
  rom[04821] = 16'hffff;
  rom[04822] = 16'hffff;
  rom[04823] = 16'hffff;
  rom[04824] = 16'hffff;
  rom[04825] = 16'hffff;
  rom[04826] = 16'hffff;
  rom[04827] = 16'hffff;
  rom[04828] = 16'hffff;
  rom[04829] = 16'hffff;
  rom[04830] = 16'hffff;
  rom[04831] = 16'hffff;
  rom[04832] = 16'hffff;
  rom[04833] = 16'hffff;
  rom[04834] = 16'hffff;
  rom[04835] = 16'hffff;
  rom[04836] = 16'hffff;
  rom[04837] = 16'hffff;
  rom[04838] = 16'hffff;
  rom[04839] = 16'hffff;
  rom[04840] = 16'hffff;
  rom[04841] = 16'hffff;
  rom[04842] = 16'hffff;
  rom[04843] = 16'hffff;
  rom[04844] = 16'hffff;
  rom[04845] = 16'hffff;
  rom[04846] = 16'hffff;
  rom[04847] = 16'hffff;
  rom[04848] = 16'hffff;
  rom[04849] = 16'hffff;
  rom[04850] = 16'hffff;
  rom[04851] = 16'hffff;
  rom[04852] = 16'hffff;
  rom[04853] = 16'hdebb;
  rom[04854] = 16'h41e7;
  rom[04855] = 16'h10a2;
  rom[04856] = 16'h10a2;
  rom[04857] = 16'h10a2;
  rom[04858] = 16'h10a3;
  rom[04859] = 16'h18a3;
  rom[04860] = 16'h10a3;
  rom[04861] = 16'h18c3;
  rom[04862] = 16'h10c2;
  rom[04863] = 16'h10c2;
  rom[04864] = 16'h08a1;
  rom[04865] = 16'h10a2;
  rom[04866] = 16'h18c3;
  rom[04867] = 16'h526b;
  rom[04868] = 16'hef5d;
  rom[04869] = 16'hfffe;
  rom[04870] = 16'hb551;
  rom[04871] = 16'hb4ac;
  rom[04872] = 16'hd58c;
  rom[04873] = 16'hf62d;
  rom[04874] = 16'hd507;
  rom[04875] = 16'hf5c9;
  rom[04876] = 16'hf586;
  rom[04877] = 16'hfda8;
  rom[04878] = 16'hf548;
  rom[04879] = 16'hf569;
  rom[04880] = 16'hf589;
  rom[04881] = 16'hfda8;
  rom[04882] = 16'hfd88;
  rom[04883] = 16'hfda8;
  rom[04884] = 16'hf587;
  rom[04885] = 16'hfda8;
  rom[04886] = 16'hfd88;
  rom[04887] = 16'hfda8;
  rom[04888] = 16'hf588;
  rom[04889] = 16'hfda8;
  rom[04890] = 16'hfd88;
  rom[04891] = 16'hfda8;
  rom[04892] = 16'hf588;
  rom[04893] = 16'hfda8;
  rom[04894] = 16'hfd88;
  rom[04895] = 16'hfda8;
  rom[04896] = 16'hf588;
  rom[04897] = 16'hfda8;
  rom[04898] = 16'hfd88;
  rom[04899] = 16'hfda8;
  rom[04900] = 16'hf588;
  rom[04901] = 16'hfda8;
  rom[04902] = 16'hfd88;
  rom[04903] = 16'hfda8;
  rom[04904] = 16'hf588;
  rom[04905] = 16'hfda8;
  rom[04906] = 16'hfd88;
  rom[04907] = 16'hfda8;
  rom[04908] = 16'hf588;
  rom[04909] = 16'hfda8;
  rom[04910] = 16'hf588;
  rom[04911] = 16'hfda8;
  rom[04912] = 16'hf588;
  rom[04913] = 16'hf5a8;
  rom[04914] = 16'hfd68;
  rom[04915] = 16'hfd88;
  rom[04916] = 16'hf568;
  rom[04917] = 16'hfd88;
  rom[04918] = 16'hf588;
  rom[04919] = 16'hfd88;
  rom[04920] = 16'hfd68;
  rom[04921] = 16'hfd48;
  rom[04922] = 16'hfd69;
  rom[04923] = 16'hfd69;
  rom[04924] = 16'hed69;
  rom[04925] = 16'hd50c;
  rom[04926] = 16'h51c4;
  rom[04927] = 16'h1882;
  rom[04928] = 16'h18a2;
  rom[04929] = 16'h18a2;
  rom[04930] = 16'h10a2;
  rom[04931] = 16'h10c2;
  rom[04932] = 16'h10a2;
  rom[04933] = 16'h10a3;
  rom[04934] = 16'h10a3;
  rom[04935] = 16'h10a2;
  rom[04936] = 16'h1081;
  rom[04937] = 16'h18c2;
  rom[04938] = 16'h1062;
  rom[04939] = 16'h18c3;
  rom[04940] = 16'h9492;
  rom[04941] = 16'hffff;
  rom[04942] = 16'hffff;
  rom[04943] = 16'hffff;
  rom[04944] = 16'hffff;
  rom[04945] = 16'hffff;
  rom[04946] = 16'hffff;
  rom[04947] = 16'hffff;
  rom[04948] = 16'hffff;
  rom[04949] = 16'hffff;
  rom[04950] = 16'hffff;
  rom[04951] = 16'hffff;
  rom[04952] = 16'hffff;
  rom[04953] = 16'hffff;
  rom[04954] = 16'hffff;
  rom[04955] = 16'hffff;
  rom[04956] = 16'hffff;
  rom[04957] = 16'hffff;
  rom[04958] = 16'hffff;
  rom[04959] = 16'hffff;
  rom[04960] = 16'hffff;
  rom[04961] = 16'hffff;
  rom[04962] = 16'hffff;
  rom[04963] = 16'hffff;
  rom[04964] = 16'hffff;
  rom[04965] = 16'hffff;
  rom[04966] = 16'hffff;
  rom[04967] = 16'hffff;
  rom[04968] = 16'hffff;
  rom[04969] = 16'hffff;
  rom[04970] = 16'hffff;
  rom[04971] = 16'hffff;
  rom[04972] = 16'hffff;
  rom[04973] = 16'hffff;
  rom[04974] = 16'hffff;
  rom[04975] = 16'hffff;
  rom[04976] = 16'hffff;
  rom[04977] = 16'hffff;
  rom[04978] = 16'hffff;
  rom[04979] = 16'hffff;
  rom[04980] = 16'hffff;
  rom[04981] = 16'hffff;
  rom[04982] = 16'hffff;
  rom[04983] = 16'hffff;
  rom[04984] = 16'hffff;
  rom[04985] = 16'hffff;
  rom[04986] = 16'hffff;
  rom[04987] = 16'hffff;
  rom[04988] = 16'hffff;
  rom[04989] = 16'hffff;
  rom[04990] = 16'hffff;
  rom[04991] = 16'hffff;
  rom[04992] = 16'hffff;
  rom[04993] = 16'hffff;
  rom[04994] = 16'hffff;
  rom[04995] = 16'hffff;
  rom[04996] = 16'hffff;
  rom[04997] = 16'hffff;
  rom[04998] = 16'hffff;
  rom[04999] = 16'hffff;
  rom[05000] = 16'hffff;
  rom[05001] = 16'hffff;
  rom[05002] = 16'hffff;
  rom[05003] = 16'hffff;
  rom[05004] = 16'hffff;
  rom[05005] = 16'hffff;
  rom[05006] = 16'hffff;
  rom[05007] = 16'hffff;
  rom[05008] = 16'hffff;
  rom[05009] = 16'hffff;
  rom[05010] = 16'hffff;
  rom[05011] = 16'hffff;
  rom[05012] = 16'hffff;
  rom[05013] = 16'hffff;
  rom[05014] = 16'hffff;
  rom[05015] = 16'hffff;
  rom[05016] = 16'hffff;
  rom[05017] = 16'hffff;
  rom[05018] = 16'hffff;
  rom[05019] = 16'hffff;
  rom[05020] = 16'hffff;
  rom[05021] = 16'hffff;
  rom[05022] = 16'hffff;
  rom[05023] = 16'hffff;
  rom[05024] = 16'hffff;
  rom[05025] = 16'hffff;
  rom[05026] = 16'hffff;
  rom[05027] = 16'hffff;
  rom[05028] = 16'hffff;
  rom[05029] = 16'hffff;
  rom[05030] = 16'hffff;
  rom[05031] = 16'hffff;
  rom[05032] = 16'hffff;
  rom[05033] = 16'hffff;
  rom[05034] = 16'hffff;
  rom[05035] = 16'hffff;
  rom[05036] = 16'hffff;
  rom[05037] = 16'hffff;
  rom[05038] = 16'hffff;
  rom[05039] = 16'hffff;
  rom[05040] = 16'hffff;
  rom[05041] = 16'hffff;
  rom[05042] = 16'hffff;
  rom[05043] = 16'hffff;
  rom[05044] = 16'hffff;
  rom[05045] = 16'hffff;
  rom[05046] = 16'hffff;
  rom[05047] = 16'hffff;
  rom[05048] = 16'hffff;
  rom[05049] = 16'hffff;
  rom[05050] = 16'hffff;
  rom[05051] = 16'hffff;
  rom[05052] = 16'hffff;
  rom[05053] = 16'he6fc;
  rom[05054] = 16'h4a49;
  rom[05055] = 16'h10a2;
  rom[05056] = 16'h18c3;
  rom[05057] = 16'h10a3;
  rom[05058] = 16'h18a3;
  rom[05059] = 16'h18a3;
  rom[05060] = 16'h10a3;
  rom[05061] = 16'h10a2;
  rom[05062] = 16'h10c2;
  rom[05063] = 16'h10c2;
  rom[05064] = 16'h08a1;
  rom[05065] = 16'h10c3;
  rom[05066] = 16'h20e5;
  rom[05067] = 16'h4a2a;
  rom[05068] = 16'hf79f;
  rom[05069] = 16'hffdd;
  rom[05070] = 16'ha44c;
  rom[05071] = 16'hac89;
  rom[05072] = 16'he5eb;
  rom[05073] = 16'hedc9;
  rom[05074] = 16'hf5a8;
  rom[05075] = 16'hf5a7;
  rom[05076] = 16'hfda6;
  rom[05077] = 16'hfd67;
  rom[05078] = 16'hfd6a;
  rom[05079] = 16'hfd69;
  rom[05080] = 16'hfd89;
  rom[05081] = 16'hfd68;
  rom[05082] = 16'hfd88;
  rom[05083] = 16'hfd88;
  rom[05084] = 16'hfdc9;
  rom[05085] = 16'hfd88;
  rom[05086] = 16'hfda9;
  rom[05087] = 16'hfd88;
  rom[05088] = 16'hfda9;
  rom[05089] = 16'hfd88;
  rom[05090] = 16'hfda9;
  rom[05091] = 16'hfda8;
  rom[05092] = 16'hfdc9;
  rom[05093] = 16'hfd88;
  rom[05094] = 16'hfda9;
  rom[05095] = 16'hfd88;
  rom[05096] = 16'hfda9;
  rom[05097] = 16'hfd88;
  rom[05098] = 16'hfda9;
  rom[05099] = 16'hfd88;
  rom[05100] = 16'hfda9;
  rom[05101] = 16'hfd88;
  rom[05102] = 16'hfda9;
  rom[05103] = 16'hfd88;
  rom[05104] = 16'hfda9;
  rom[05105] = 16'hfd88;
  rom[05106] = 16'hfda9;
  rom[05107] = 16'hfd88;
  rom[05108] = 16'hfda9;
  rom[05109] = 16'hfd88;
  rom[05110] = 16'hfda9;
  rom[05111] = 16'hfd88;
  rom[05112] = 16'hfda9;
  rom[05113] = 16'hfd88;
  rom[05114] = 16'hfd88;
  rom[05115] = 16'hfd68;
  rom[05116] = 16'hfd88;
  rom[05117] = 16'hfd88;
  rom[05118] = 16'hf589;
  rom[05119] = 16'hf568;
  rom[05120] = 16'hfd89;
  rom[05121] = 16'hfd48;
  rom[05122] = 16'hfd8a;
  rom[05123] = 16'hfd49;
  rom[05124] = 16'hfd8a;
  rom[05125] = 16'hc4aa;
  rom[05126] = 16'h51e4;
  rom[05127] = 16'h20a1;
  rom[05128] = 16'h1882;
  rom[05129] = 16'h18c2;
  rom[05130] = 16'h10c3;
  rom[05131] = 16'h10c2;
  rom[05132] = 16'h10c3;
  rom[05133] = 16'h10a3;
  rom[05134] = 16'h10c3;
  rom[05135] = 16'h10a2;
  rom[05136] = 16'h18e3;
  rom[05137] = 16'h10a2;
  rom[05138] = 16'h18c3;
  rom[05139] = 16'h2945;
  rom[05140] = 16'hb576;
  rom[05141] = 16'hffff;
  rom[05142] = 16'hffff;
  rom[05143] = 16'hffff;
  rom[05144] = 16'hffff;
  rom[05145] = 16'hffff;
  rom[05146] = 16'hffff;
  rom[05147] = 16'hffff;
  rom[05148] = 16'hffff;
  rom[05149] = 16'hffff;
  rom[05150] = 16'hffff;
  rom[05151] = 16'hffff;
  rom[05152] = 16'hffff;
  rom[05153] = 16'hffff;
  rom[05154] = 16'hffff;
  rom[05155] = 16'hffff;
  rom[05156] = 16'hffff;
  rom[05157] = 16'hffff;
  rom[05158] = 16'hffff;
  rom[05159] = 16'hffff;
  rom[05160] = 16'hffff;
  rom[05161] = 16'hffff;
  rom[05162] = 16'hffff;
  rom[05163] = 16'hffff;
  rom[05164] = 16'hffff;
  rom[05165] = 16'hffff;
  rom[05166] = 16'hffff;
  rom[05167] = 16'hffff;
  rom[05168] = 16'hffff;
  rom[05169] = 16'hffff;
  rom[05170] = 16'hffff;
  rom[05171] = 16'hffff;
  rom[05172] = 16'hffff;
  rom[05173] = 16'hffff;
  rom[05174] = 16'hffff;
  rom[05175] = 16'hffff;
  rom[05176] = 16'hffff;
  rom[05177] = 16'hffff;
  rom[05178] = 16'hffff;
  rom[05179] = 16'hffff;
  rom[05180] = 16'hffff;
  rom[05181] = 16'hffff;
  rom[05182] = 16'hffff;
  rom[05183] = 16'hffff;
  rom[05184] = 16'hffff;
  rom[05185] = 16'hffff;
  rom[05186] = 16'hffff;
  rom[05187] = 16'hffff;
  rom[05188] = 16'hffff;
  rom[05189] = 16'hffff;
  rom[05190] = 16'hffff;
  rom[05191] = 16'hffff;
  rom[05192] = 16'hffff;
  rom[05193] = 16'hffff;
  rom[05194] = 16'hffff;
  rom[05195] = 16'hffff;
  rom[05196] = 16'hffff;
  rom[05197] = 16'hffff;
  rom[05198] = 16'hffff;
  rom[05199] = 16'hffff;
  rom[05200] = 16'hffff;
  rom[05201] = 16'hffff;
  rom[05202] = 16'hffff;
  rom[05203] = 16'hffff;
  rom[05204] = 16'hffff;
  rom[05205] = 16'hffff;
  rom[05206] = 16'hffff;
  rom[05207] = 16'hffff;
  rom[05208] = 16'hffff;
  rom[05209] = 16'hffff;
  rom[05210] = 16'hffff;
  rom[05211] = 16'hffff;
  rom[05212] = 16'hffff;
  rom[05213] = 16'hffff;
  rom[05214] = 16'hffff;
  rom[05215] = 16'hffff;
  rom[05216] = 16'hffff;
  rom[05217] = 16'hffff;
  rom[05218] = 16'hffff;
  rom[05219] = 16'hffff;
  rom[05220] = 16'hffff;
  rom[05221] = 16'hffff;
  rom[05222] = 16'hffff;
  rom[05223] = 16'hffff;
  rom[05224] = 16'hffff;
  rom[05225] = 16'hffff;
  rom[05226] = 16'hffff;
  rom[05227] = 16'hffff;
  rom[05228] = 16'hffff;
  rom[05229] = 16'hffff;
  rom[05230] = 16'hffff;
  rom[05231] = 16'hffff;
  rom[05232] = 16'hffff;
  rom[05233] = 16'hffff;
  rom[05234] = 16'hffff;
  rom[05235] = 16'hffff;
  rom[05236] = 16'hffff;
  rom[05237] = 16'hffff;
  rom[05238] = 16'hffff;
  rom[05239] = 16'hffff;
  rom[05240] = 16'hffff;
  rom[05241] = 16'hffff;
  rom[05242] = 16'hffff;
  rom[05243] = 16'hffff;
  rom[05244] = 16'hffff;
  rom[05245] = 16'hffff;
  rom[05246] = 16'hffff;
  rom[05247] = 16'hffff;
  rom[05248] = 16'hffff;
  rom[05249] = 16'hffff;
  rom[05250] = 16'hffff;
  rom[05251] = 16'hffff;
  rom[05252] = 16'hffff;
  rom[05253] = 16'hf79e;
  rom[05254] = 16'h4a69;
  rom[05255] = 16'h10a2;
  rom[05256] = 16'h10a2;
  rom[05257] = 16'h10a2;
  rom[05258] = 16'h18a3;
  rom[05259] = 16'h18a3;
  rom[05260] = 16'h18a2;
  rom[05261] = 16'h18c2;
  rom[05262] = 16'h10e2;
  rom[05263] = 16'h10a2;
  rom[05264] = 16'h08a1;
  rom[05265] = 16'h10c3;
  rom[05266] = 16'h10c3;
  rom[05267] = 16'h524a;
  rom[05268] = 16'hef3c;
  rom[05269] = 16'hde56;
  rom[05270] = 16'h7b05;
  rom[05271] = 16'hcd2b;
  rom[05272] = 16'hee0a;
  rom[05273] = 16'heda8;
  rom[05274] = 16'heda7;
  rom[05275] = 16'hf5a7;
  rom[05276] = 16'hfda6;
  rom[05277] = 16'hfda8;
  rom[05278] = 16'hfd69;
  rom[05279] = 16'hfd89;
  rom[05280] = 16'hfd68;
  rom[05281] = 16'hfda8;
  rom[05282] = 16'hf588;
  rom[05283] = 16'hf5a7;
  rom[05284] = 16'hfd88;
  rom[05285] = 16'hfda8;
  rom[05286] = 16'hf588;
  rom[05287] = 16'hfda8;
  rom[05288] = 16'hfd88;
  rom[05289] = 16'hfda8;
  rom[05290] = 16'hf5a8;
  rom[05291] = 16'hfdc8;
  rom[05292] = 16'hfda8;
  rom[05293] = 16'hfdc8;
  rom[05294] = 16'hf5a8;
  rom[05295] = 16'hfda8;
  rom[05296] = 16'hfda9;
  rom[05297] = 16'hfdc9;
  rom[05298] = 16'hf5a9;
  rom[05299] = 16'hfdc8;
  rom[05300] = 16'hfda8;
  rom[05301] = 16'hfda8;
  rom[05302] = 16'hf588;
  rom[05303] = 16'hfda8;
  rom[05304] = 16'hfd88;
  rom[05305] = 16'hfda8;
  rom[05306] = 16'hf5a8;
  rom[05307] = 16'hfda8;
  rom[05308] = 16'hfd88;
  rom[05309] = 16'hfda8;
  rom[05310] = 16'hf588;
  rom[05311] = 16'hfda8;
  rom[05312] = 16'hfd88;
  rom[05313] = 16'hfda8;
  rom[05314] = 16'hf587;
  rom[05315] = 16'hfd87;
  rom[05316] = 16'hfd87;
  rom[05317] = 16'hfda8;
  rom[05318] = 16'hed88;
  rom[05319] = 16'hf588;
  rom[05320] = 16'hfd49;
  rom[05321] = 16'hfd49;
  rom[05322] = 16'hfd69;
  rom[05323] = 16'hfd49;
  rom[05324] = 16'hf589;
  rom[05325] = 16'hbc69;
  rom[05326] = 16'h3921;
  rom[05327] = 16'h1881;
  rom[05328] = 16'h18a2;
  rom[05329] = 16'h18c3;
  rom[05330] = 16'h10a2;
  rom[05331] = 16'h10c3;
  rom[05332] = 16'h10a3;
  rom[05333] = 16'h10a3;
  rom[05334] = 16'h10a2;
  rom[05335] = 16'h10e3;
  rom[05336] = 16'h10c2;
  rom[05337] = 16'h18c3;
  rom[05338] = 16'h10a2;
  rom[05339] = 16'h39e7;
  rom[05340] = 16'hbdf8;
  rom[05341] = 16'hffff;
  rom[05342] = 16'hffff;
  rom[05343] = 16'hffff;
  rom[05344] = 16'hffff;
  rom[05345] = 16'hffff;
  rom[05346] = 16'hffff;
  rom[05347] = 16'hffff;
  rom[05348] = 16'hffff;
  rom[05349] = 16'hffff;
  rom[05350] = 16'hffff;
  rom[05351] = 16'hffff;
  rom[05352] = 16'hffff;
  rom[05353] = 16'hffff;
  rom[05354] = 16'hffff;
  rom[05355] = 16'hffff;
  rom[05356] = 16'hffff;
  rom[05357] = 16'hffff;
  rom[05358] = 16'hffff;
  rom[05359] = 16'hffff;
  rom[05360] = 16'hffff;
  rom[05361] = 16'hffff;
  rom[05362] = 16'hffff;
  rom[05363] = 16'hffff;
  rom[05364] = 16'hffff;
  rom[05365] = 16'hffff;
  rom[05366] = 16'hffff;
  rom[05367] = 16'hffff;
  rom[05368] = 16'hffff;
  rom[05369] = 16'hffff;
  rom[05370] = 16'hffff;
  rom[05371] = 16'hffff;
  rom[05372] = 16'hffff;
  rom[05373] = 16'hffff;
  rom[05374] = 16'hffff;
  rom[05375] = 16'hffff;
  rom[05376] = 16'hffff;
  rom[05377] = 16'hffff;
  rom[05378] = 16'hffff;
  rom[05379] = 16'hffff;
  rom[05380] = 16'hffff;
  rom[05381] = 16'hffff;
  rom[05382] = 16'hffff;
  rom[05383] = 16'hffff;
  rom[05384] = 16'hffff;
  rom[05385] = 16'hffff;
  rom[05386] = 16'hffff;
  rom[05387] = 16'hffff;
  rom[05388] = 16'hffff;
  rom[05389] = 16'hffff;
  rom[05390] = 16'hffff;
  rom[05391] = 16'hffff;
  rom[05392] = 16'hffff;
  rom[05393] = 16'hffff;
  rom[05394] = 16'hffff;
  rom[05395] = 16'hffff;
  rom[05396] = 16'hffff;
  rom[05397] = 16'hffff;
  rom[05398] = 16'hffff;
  rom[05399] = 16'hffff;
  rom[05400] = 16'hffff;
  rom[05401] = 16'hffff;
  rom[05402] = 16'hffff;
  rom[05403] = 16'hffff;
  rom[05404] = 16'hffff;
  rom[05405] = 16'hffff;
  rom[05406] = 16'hffff;
  rom[05407] = 16'hffff;
  rom[05408] = 16'hffff;
  rom[05409] = 16'hffff;
  rom[05410] = 16'hffff;
  rom[05411] = 16'hffff;
  rom[05412] = 16'hffff;
  rom[05413] = 16'hffff;
  rom[05414] = 16'hffff;
  rom[05415] = 16'hffff;
  rom[05416] = 16'hffff;
  rom[05417] = 16'hffff;
  rom[05418] = 16'hffff;
  rom[05419] = 16'hffff;
  rom[05420] = 16'hffff;
  rom[05421] = 16'hffff;
  rom[05422] = 16'hffff;
  rom[05423] = 16'hffff;
  rom[05424] = 16'hffff;
  rom[05425] = 16'hffff;
  rom[05426] = 16'hffff;
  rom[05427] = 16'hffff;
  rom[05428] = 16'hffff;
  rom[05429] = 16'hffff;
  rom[05430] = 16'hffff;
  rom[05431] = 16'hffff;
  rom[05432] = 16'hffff;
  rom[05433] = 16'hffff;
  rom[05434] = 16'hffff;
  rom[05435] = 16'hffff;
  rom[05436] = 16'hffff;
  rom[05437] = 16'hffff;
  rom[05438] = 16'hffff;
  rom[05439] = 16'hffff;
  rom[05440] = 16'hffff;
  rom[05441] = 16'hffff;
  rom[05442] = 16'hffff;
  rom[05443] = 16'hffff;
  rom[05444] = 16'hffff;
  rom[05445] = 16'hffff;
  rom[05446] = 16'hffff;
  rom[05447] = 16'hffff;
  rom[05448] = 16'hffff;
  rom[05449] = 16'hffff;
  rom[05450] = 16'hffff;
  rom[05451] = 16'hffff;
  rom[05452] = 16'hffff;
  rom[05453] = 16'hffdf;
  rom[05454] = 16'h738e;
  rom[05455] = 16'h18e3;
  rom[05456] = 16'h10c2;
  rom[05457] = 16'h10a2;
  rom[05458] = 16'h18c3;
  rom[05459] = 16'h18a3;
  rom[05460] = 16'h18a3;
  rom[05461] = 16'h18a2;
  rom[05462] = 16'h18c3;
  rom[05463] = 16'h10a2;
  rom[05464] = 16'h10a2;
  rom[05465] = 16'h18c3;
  rom[05466] = 16'h1082;
  rom[05467] = 16'h4a07;
  rom[05468] = 16'hacb1;
  rom[05469] = 16'h7b27;
  rom[05470] = 16'hac28;
  rom[05471] = 16'he56b;
  rom[05472] = 16'hf5aa;
  rom[05473] = 16'hf589;
  rom[05474] = 16'hfda9;
  rom[05475] = 16'hfda8;
  rom[05476] = 16'hfda7;
  rom[05477] = 16'hf587;
  rom[05478] = 16'hfd89;
  rom[05479] = 16'hfd69;
  rom[05480] = 16'hfd89;
  rom[05481] = 16'hfd88;
  rom[05482] = 16'hfda8;
  rom[05483] = 16'hfda8;
  rom[05484] = 16'hfda9;
  rom[05485] = 16'hfda8;
  rom[05486] = 16'hfda9;
  rom[05487] = 16'hfda9;
  rom[05488] = 16'hfda9;
  rom[05489] = 16'hfd88;
  rom[05490] = 16'hfdc9;
  rom[05491] = 16'hfda8;
  rom[05492] = 16'hfdc9;
  rom[05493] = 16'hfda8;
  rom[05494] = 16'hfdc9;
  rom[05495] = 16'hfda9;
  rom[05496] = 16'hfdca;
  rom[05497] = 16'hfda8;
  rom[05498] = 16'hfdc9;
  rom[05499] = 16'hfda8;
  rom[05500] = 16'hfdc9;
  rom[05501] = 16'hfda8;
  rom[05502] = 16'hfdc9;
  rom[05503] = 16'hfda8;
  rom[05504] = 16'hfdc9;
  rom[05505] = 16'hfda8;
  rom[05506] = 16'hfdc9;
  rom[05507] = 16'hfda8;
  rom[05508] = 16'hfdc9;
  rom[05509] = 16'hfda8;
  rom[05510] = 16'hfdc9;
  rom[05511] = 16'hfda8;
  rom[05512] = 16'hfda9;
  rom[05513] = 16'hfd88;
  rom[05514] = 16'hfda9;
  rom[05515] = 16'hfd87;
  rom[05516] = 16'hfda8;
  rom[05517] = 16'hf5a7;
  rom[05518] = 16'hf5a9;
  rom[05519] = 16'hfd88;
  rom[05520] = 16'hfd69;
  rom[05521] = 16'hfd69;
  rom[05522] = 16'hfd69;
  rom[05523] = 16'hf568;
  rom[05524] = 16'hf5aa;
  rom[05525] = 16'hac28;
  rom[05526] = 16'h3101;
  rom[05527] = 16'h18a1;
  rom[05528] = 16'h20a2;
  rom[05529] = 16'h18a2;
  rom[05530] = 16'h10c3;
  rom[05531] = 16'h10c3;
  rom[05532] = 16'h18c3;
  rom[05533] = 16'h10a3;
  rom[05534] = 16'h10c2;
  rom[05535] = 16'h10c2;
  rom[05536] = 16'h18c3;
  rom[05537] = 16'h10c2;
  rom[05538] = 16'h10a2;
  rom[05539] = 16'h39e7;
  rom[05540] = 16'hdebb;
  rom[05541] = 16'hffff;
  rom[05542] = 16'hffff;
  rom[05543] = 16'hffff;
  rom[05544] = 16'hffff;
  rom[05545] = 16'hffff;
  rom[05546] = 16'hffff;
  rom[05547] = 16'hffff;
  rom[05548] = 16'hffff;
  rom[05549] = 16'hffff;
  rom[05550] = 16'hffff;
  rom[05551] = 16'hffff;
  rom[05552] = 16'hffff;
  rom[05553] = 16'hffff;
  rom[05554] = 16'hffff;
  rom[05555] = 16'hffff;
  rom[05556] = 16'hffff;
  rom[05557] = 16'hffff;
  rom[05558] = 16'hffff;
  rom[05559] = 16'hffff;
  rom[05560] = 16'hffff;
  rom[05561] = 16'hffff;
  rom[05562] = 16'hffff;
  rom[05563] = 16'hffff;
  rom[05564] = 16'hffff;
  rom[05565] = 16'hffff;
  rom[05566] = 16'hffff;
  rom[05567] = 16'hffff;
  rom[05568] = 16'hffff;
  rom[05569] = 16'hffff;
  rom[05570] = 16'hffff;
  rom[05571] = 16'hffff;
  rom[05572] = 16'hffff;
  rom[05573] = 16'hffff;
  rom[05574] = 16'hffff;
  rom[05575] = 16'hffff;
  rom[05576] = 16'hffff;
  rom[05577] = 16'hffff;
  rom[05578] = 16'hffff;
  rom[05579] = 16'hffff;
  rom[05580] = 16'hffff;
  rom[05581] = 16'hffff;
  rom[05582] = 16'hffff;
  rom[05583] = 16'hffff;
  rom[05584] = 16'hffff;
  rom[05585] = 16'hffff;
  rom[05586] = 16'hffff;
  rom[05587] = 16'hffff;
  rom[05588] = 16'hffff;
  rom[05589] = 16'hffff;
  rom[05590] = 16'hffff;
  rom[05591] = 16'hffff;
  rom[05592] = 16'hffff;
  rom[05593] = 16'hffff;
  rom[05594] = 16'hffff;
  rom[05595] = 16'hffff;
  rom[05596] = 16'hffff;
  rom[05597] = 16'hffff;
  rom[05598] = 16'hffff;
  rom[05599] = 16'hffff;
  rom[05600] = 16'hffff;
  rom[05601] = 16'hffff;
  rom[05602] = 16'hffff;
  rom[05603] = 16'hffff;
  rom[05604] = 16'hffff;
  rom[05605] = 16'hffff;
  rom[05606] = 16'hffff;
  rom[05607] = 16'hffff;
  rom[05608] = 16'hffff;
  rom[05609] = 16'hffff;
  rom[05610] = 16'hffff;
  rom[05611] = 16'hffff;
  rom[05612] = 16'hffff;
  rom[05613] = 16'hffff;
  rom[05614] = 16'hffff;
  rom[05615] = 16'hffff;
  rom[05616] = 16'hffff;
  rom[05617] = 16'hffff;
  rom[05618] = 16'hffff;
  rom[05619] = 16'hffff;
  rom[05620] = 16'hffff;
  rom[05621] = 16'hffff;
  rom[05622] = 16'hffff;
  rom[05623] = 16'hffff;
  rom[05624] = 16'hffff;
  rom[05625] = 16'hffff;
  rom[05626] = 16'hffff;
  rom[05627] = 16'hffff;
  rom[05628] = 16'hffff;
  rom[05629] = 16'hffff;
  rom[05630] = 16'hffff;
  rom[05631] = 16'hffff;
  rom[05632] = 16'hffff;
  rom[05633] = 16'hffff;
  rom[05634] = 16'hffff;
  rom[05635] = 16'hffff;
  rom[05636] = 16'hffff;
  rom[05637] = 16'hffff;
  rom[05638] = 16'hffff;
  rom[05639] = 16'hffff;
  rom[05640] = 16'hffff;
  rom[05641] = 16'hffff;
  rom[05642] = 16'hffff;
  rom[05643] = 16'hffff;
  rom[05644] = 16'hffff;
  rom[05645] = 16'hffff;
  rom[05646] = 16'hffff;
  rom[05647] = 16'hffff;
  rom[05648] = 16'hffff;
  rom[05649] = 16'hffff;
  rom[05650] = 16'hffff;
  rom[05651] = 16'hffff;
  rom[05652] = 16'hffdf;
  rom[05653] = 16'hffff;
  rom[05654] = 16'h94b2;
  rom[05655] = 16'h18e3;
  rom[05656] = 16'h10a1;
  rom[05657] = 16'h10c1;
  rom[05658] = 16'h18a2;
  rom[05659] = 16'h18a2;
  rom[05660] = 16'h18a3;
  rom[05661] = 16'h18a3;
  rom[05662] = 16'h1084;
  rom[05663] = 16'h18c4;
  rom[05664] = 16'h0861;
  rom[05665] = 16'h18a2;
  rom[05666] = 16'h1881;
  rom[05667] = 16'h30e2;
  rom[05668] = 16'h6aa7;
  rom[05669] = 16'hbccc;
  rom[05670] = 16'he58c;
  rom[05671] = 16'hed4a;
  rom[05672] = 16'hfdaa;
  rom[05673] = 16'hfd69;
  rom[05674] = 16'hfda9;
  rom[05675] = 16'hfd89;
  rom[05676] = 16'hf5a8;
  rom[05677] = 16'hfda8;
  rom[05678] = 16'hfda9;
  rom[05679] = 16'hfd89;
  rom[05680] = 16'hf588;
  rom[05681] = 16'hfd88;
  rom[05682] = 16'hf5a8;
  rom[05683] = 16'hfdc8;
  rom[05684] = 16'hf5a8;
  rom[05685] = 16'hfdc9;
  rom[05686] = 16'hfda9;
  rom[05687] = 16'hfdc9;
  rom[05688] = 16'hf5a9;
  rom[05689] = 16'hfda8;
  rom[05690] = 16'hfda8;
  rom[05691] = 16'hfdc8;
  rom[05692] = 16'hf5a8;
  rom[05693] = 16'hfdc9;
  rom[05694] = 16'hfda8;
  rom[05695] = 16'hfdc9;
  rom[05696] = 16'hf5a9;
  rom[05697] = 16'hfdc9;
  rom[05698] = 16'hfda8;
  rom[05699] = 16'hfdc8;
  rom[05700] = 16'hf5a8;
  rom[05701] = 16'hfdc8;
  rom[05702] = 16'hfda8;
  rom[05703] = 16'hfdc8;
  rom[05704] = 16'hf5a8;
  rom[05705] = 16'hfdc8;
  rom[05706] = 16'hfda8;
  rom[05707] = 16'hfdc8;
  rom[05708] = 16'hf5a8;
  rom[05709] = 16'hfdc8;
  rom[05710] = 16'hfda8;
  rom[05711] = 16'hfdc8;
  rom[05712] = 16'hf588;
  rom[05713] = 16'hfda9;
  rom[05714] = 16'hfd68;
  rom[05715] = 16'hfda8;
  rom[05716] = 16'hf5a7;
  rom[05717] = 16'hf5c7;
  rom[05718] = 16'hf5a8;
  rom[05719] = 16'hfda9;
  rom[05720] = 16'hf568;
  rom[05721] = 16'hfd69;
  rom[05722] = 16'hfd68;
  rom[05723] = 16'hf589;
  rom[05724] = 16'he569;
  rom[05725] = 16'h9bc7;
  rom[05726] = 16'h28e0;
  rom[05727] = 16'h20c1;
  rom[05728] = 16'h18a1;
  rom[05729] = 16'h18a2;
  rom[05730] = 16'h10a3;
  rom[05731] = 16'h10c3;
  rom[05732] = 16'h10a3;
  rom[05733] = 16'h10a3;
  rom[05734] = 16'h10a2;
  rom[05735] = 16'h10c3;
  rom[05736] = 16'h10a2;
  rom[05737] = 16'h10c3;
  rom[05738] = 16'h10c2;
  rom[05739] = 16'h4a49;
  rom[05740] = 16'he73c;
  rom[05741] = 16'hffff;
  rom[05742] = 16'hffff;
  rom[05743] = 16'hffff;
  rom[05744] = 16'hffff;
  rom[05745] = 16'hffff;
  rom[05746] = 16'hffff;
  rom[05747] = 16'hffff;
  rom[05748] = 16'hffff;
  rom[05749] = 16'hffff;
  rom[05750] = 16'hffff;
  rom[05751] = 16'hffff;
  rom[05752] = 16'hffff;
  rom[05753] = 16'hffff;
  rom[05754] = 16'hffff;
  rom[05755] = 16'hffff;
  rom[05756] = 16'hffff;
  rom[05757] = 16'hffff;
  rom[05758] = 16'hffff;
  rom[05759] = 16'hffff;
  rom[05760] = 16'hffff;
  rom[05761] = 16'hffff;
  rom[05762] = 16'hffff;
  rom[05763] = 16'hffff;
  rom[05764] = 16'hffff;
  rom[05765] = 16'hffff;
  rom[05766] = 16'hffff;
  rom[05767] = 16'hffff;
  rom[05768] = 16'hffff;
  rom[05769] = 16'hffff;
  rom[05770] = 16'hffff;
  rom[05771] = 16'hffff;
  rom[05772] = 16'hffff;
  rom[05773] = 16'hffff;
  rom[05774] = 16'hffff;
  rom[05775] = 16'hffff;
  rom[05776] = 16'hffff;
  rom[05777] = 16'hffff;
  rom[05778] = 16'hffff;
  rom[05779] = 16'hffff;
  rom[05780] = 16'hffff;
  rom[05781] = 16'hffff;
  rom[05782] = 16'hffff;
  rom[05783] = 16'hffff;
  rom[05784] = 16'hffff;
  rom[05785] = 16'hffff;
  rom[05786] = 16'hffff;
  rom[05787] = 16'hffff;
  rom[05788] = 16'hffff;
  rom[05789] = 16'hffff;
  rom[05790] = 16'hffff;
  rom[05791] = 16'hffff;
  rom[05792] = 16'hffff;
  rom[05793] = 16'hffff;
  rom[05794] = 16'hffff;
  rom[05795] = 16'hffff;
  rom[05796] = 16'hffff;
  rom[05797] = 16'hffff;
  rom[05798] = 16'hffff;
  rom[05799] = 16'hffff;
  rom[05800] = 16'hffff;
  rom[05801] = 16'hffff;
  rom[05802] = 16'hffff;
  rom[05803] = 16'hffff;
  rom[05804] = 16'hffff;
  rom[05805] = 16'hffff;
  rom[05806] = 16'hffff;
  rom[05807] = 16'hffff;
  rom[05808] = 16'hffff;
  rom[05809] = 16'hffff;
  rom[05810] = 16'hffff;
  rom[05811] = 16'hffff;
  rom[05812] = 16'hffff;
  rom[05813] = 16'hffff;
  rom[05814] = 16'hffff;
  rom[05815] = 16'hffff;
  rom[05816] = 16'hffff;
  rom[05817] = 16'hffff;
  rom[05818] = 16'hffff;
  rom[05819] = 16'hffff;
  rom[05820] = 16'hffff;
  rom[05821] = 16'hffff;
  rom[05822] = 16'hffff;
  rom[05823] = 16'hffff;
  rom[05824] = 16'hffff;
  rom[05825] = 16'hffff;
  rom[05826] = 16'hffff;
  rom[05827] = 16'hffff;
  rom[05828] = 16'hffff;
  rom[05829] = 16'hffff;
  rom[05830] = 16'hffff;
  rom[05831] = 16'hffff;
  rom[05832] = 16'hffff;
  rom[05833] = 16'hffff;
  rom[05834] = 16'hffff;
  rom[05835] = 16'hffff;
  rom[05836] = 16'hffff;
  rom[05837] = 16'hffff;
  rom[05838] = 16'hffff;
  rom[05839] = 16'hffff;
  rom[05840] = 16'hffff;
  rom[05841] = 16'hffff;
  rom[05842] = 16'hffff;
  rom[05843] = 16'hffff;
  rom[05844] = 16'hffff;
  rom[05845] = 16'hffff;
  rom[05846] = 16'hffff;
  rom[05847] = 16'hffff;
  rom[05848] = 16'hffff;
  rom[05849] = 16'hffff;
  rom[05850] = 16'hffff;
  rom[05851] = 16'hffff;
  rom[05852] = 16'hffff;
  rom[05853] = 16'hffff;
  rom[05854] = 16'hc5f8;
  rom[05855] = 16'h18c2;
  rom[05856] = 16'h10c1;
  rom[05857] = 16'h10c1;
  rom[05858] = 16'h18c2;
  rom[05859] = 16'h18a2;
  rom[05860] = 16'h18a4;
  rom[05861] = 16'h1884;
  rom[05862] = 16'h18a5;
  rom[05863] = 16'h1884;
  rom[05864] = 16'h1883;
  rom[05865] = 16'h20a2;
  rom[05866] = 16'h28a2;
  rom[05867] = 16'h28a0;
  rom[05868] = 16'hac4c;
  rom[05869] = 16'he5ad;
  rom[05870] = 16'hf5ac;
  rom[05871] = 16'hfd89;
  rom[05872] = 16'hfda9;
  rom[05873] = 16'hfd68;
  rom[05874] = 16'hfdaa;
  rom[05875] = 16'hfd89;
  rom[05876] = 16'hfdc9;
  rom[05877] = 16'hfda8;
  rom[05878] = 16'hfda9;
  rom[05879] = 16'hfd89;
  rom[05880] = 16'hfda9;
  rom[05881] = 16'hfd88;
  rom[05882] = 16'hfda9;
  rom[05883] = 16'hfda8;
  rom[05884] = 16'hfdc9;
  rom[05885] = 16'hfda9;
  rom[05886] = 16'hfdca;
  rom[05887] = 16'hfda9;
  rom[05888] = 16'hfdca;
  rom[05889] = 16'hfda8;
  rom[05890] = 16'hfdc9;
  rom[05891] = 16'hfda8;
  rom[05892] = 16'hfdc9;
  rom[05893] = 16'hfda8;
  rom[05894] = 16'hfdc9;
  rom[05895] = 16'hfda9;
  rom[05896] = 16'hfdca;
  rom[05897] = 16'hfda8;
  rom[05898] = 16'hfdc9;
  rom[05899] = 16'hfda8;
  rom[05900] = 16'hfdc9;
  rom[05901] = 16'hfda8;
  rom[05902] = 16'hfdc9;
  rom[05903] = 16'hfda8;
  rom[05904] = 16'hfdc9;
  rom[05905] = 16'hfda8;
  rom[05906] = 16'hfdc9;
  rom[05907] = 16'hfda8;
  rom[05908] = 16'hfdc9;
  rom[05909] = 16'hfda8;
  rom[05910] = 16'hfdc9;
  rom[05911] = 16'hfda8;
  rom[05912] = 16'hfda9;
  rom[05913] = 16'hfd89;
  rom[05914] = 16'hfdaa;
  rom[05915] = 16'hfd88;
  rom[05916] = 16'hfda9;
  rom[05917] = 16'hf5a8;
  rom[05918] = 16'hf5a8;
  rom[05919] = 16'hfd88;
  rom[05920] = 16'hfd89;
  rom[05921] = 16'hfd68;
  rom[05922] = 16'hfd89;
  rom[05923] = 16'hf5ca;
  rom[05924] = 16'he56a;
  rom[05925] = 16'h8326;
  rom[05926] = 16'h3101;
  rom[05927] = 16'h18a1;
  rom[05928] = 16'h18a2;
  rom[05929] = 16'h18a2;
  rom[05930] = 16'h10a3;
  rom[05931] = 16'h10c3;
  rom[05932] = 16'h10a3;
  rom[05933] = 16'h10a3;
  rom[05934] = 16'h10c2;
  rom[05935] = 16'h10a2;
  rom[05936] = 16'h10c3;
  rom[05937] = 16'h10a2;
  rom[05938] = 16'h18e3;
  rom[05939] = 16'h738e;
  rom[05940] = 16'hffbf;
  rom[05941] = 16'hffff;
  rom[05942] = 16'hffff;
  rom[05943] = 16'hffff;
  rom[05944] = 16'hffff;
  rom[05945] = 16'hffff;
  rom[05946] = 16'hffff;
  rom[05947] = 16'hffff;
  rom[05948] = 16'hffff;
  rom[05949] = 16'hffff;
  rom[05950] = 16'hffff;
  rom[05951] = 16'hffff;
  rom[05952] = 16'hffff;
  rom[05953] = 16'hffff;
  rom[05954] = 16'hffff;
  rom[05955] = 16'hffff;
  rom[05956] = 16'hffff;
  rom[05957] = 16'hffff;
  rom[05958] = 16'hffff;
  rom[05959] = 16'hffff;
  rom[05960] = 16'hffff;
  rom[05961] = 16'hffff;
  rom[05962] = 16'hffff;
  rom[05963] = 16'hffff;
  rom[05964] = 16'hffff;
  rom[05965] = 16'hffff;
  rom[05966] = 16'hffff;
  rom[05967] = 16'hffff;
  rom[05968] = 16'hffff;
  rom[05969] = 16'hffff;
  rom[05970] = 16'hffff;
  rom[05971] = 16'hffff;
  rom[05972] = 16'hffff;
  rom[05973] = 16'hffff;
  rom[05974] = 16'hffff;
  rom[05975] = 16'hffff;
  rom[05976] = 16'hffff;
  rom[05977] = 16'hffff;
  rom[05978] = 16'hffff;
  rom[05979] = 16'hffff;
  rom[05980] = 16'hffff;
  rom[05981] = 16'hffff;
  rom[05982] = 16'hffff;
  rom[05983] = 16'hffff;
  rom[05984] = 16'hffff;
  rom[05985] = 16'hffff;
  rom[05986] = 16'hffff;
  rom[05987] = 16'hffff;
  rom[05988] = 16'hffff;
  rom[05989] = 16'hffff;
  rom[05990] = 16'hffff;
  rom[05991] = 16'hffff;
  rom[05992] = 16'hffff;
  rom[05993] = 16'hffff;
  rom[05994] = 16'hffff;
  rom[05995] = 16'hffff;
  rom[05996] = 16'hffff;
  rom[05997] = 16'hffff;
  rom[05998] = 16'hffff;
  rom[05999] = 16'hffff;
  rom[06000] = 16'hffff;
  rom[06001] = 16'hffff;
  rom[06002] = 16'hffff;
  rom[06003] = 16'hffff;
  rom[06004] = 16'hffff;
  rom[06005] = 16'hffff;
  rom[06006] = 16'hffff;
  rom[06007] = 16'hffff;
  rom[06008] = 16'hffff;
  rom[06009] = 16'hffff;
  rom[06010] = 16'hffff;
  rom[06011] = 16'hffff;
  rom[06012] = 16'hffff;
  rom[06013] = 16'hffff;
  rom[06014] = 16'hffff;
  rom[06015] = 16'hffff;
  rom[06016] = 16'hffff;
  rom[06017] = 16'hffff;
  rom[06018] = 16'hffff;
  rom[06019] = 16'hffff;
  rom[06020] = 16'hffff;
  rom[06021] = 16'hffff;
  rom[06022] = 16'hffff;
  rom[06023] = 16'hffff;
  rom[06024] = 16'hffff;
  rom[06025] = 16'hffff;
  rom[06026] = 16'hffff;
  rom[06027] = 16'hffff;
  rom[06028] = 16'hffff;
  rom[06029] = 16'hffff;
  rom[06030] = 16'hffff;
  rom[06031] = 16'hffff;
  rom[06032] = 16'hffff;
  rom[06033] = 16'hffff;
  rom[06034] = 16'hffff;
  rom[06035] = 16'hffff;
  rom[06036] = 16'hffff;
  rom[06037] = 16'hffff;
  rom[06038] = 16'hffff;
  rom[06039] = 16'hffff;
  rom[06040] = 16'hffff;
  rom[06041] = 16'hffff;
  rom[06042] = 16'hffff;
  rom[06043] = 16'hffff;
  rom[06044] = 16'hffff;
  rom[06045] = 16'hffff;
  rom[06046] = 16'hffff;
  rom[06047] = 16'hffff;
  rom[06048] = 16'hffff;
  rom[06049] = 16'hffff;
  rom[06050] = 16'hffff;
  rom[06051] = 16'hffff;
  rom[06052] = 16'hffff;
  rom[06053] = 16'hffff;
  rom[06054] = 16'hdebb;
  rom[06055] = 16'h2965;
  rom[06056] = 16'h10a1;
  rom[06057] = 16'h18e1;
  rom[06058] = 16'h10a1;
  rom[06059] = 16'h18a2;
  rom[06060] = 16'h18a3;
  rom[06061] = 16'h18a4;
  rom[06062] = 16'h1884;
  rom[06063] = 16'h18a4;
  rom[06064] = 16'h1883;
  rom[06065] = 16'h1881;
  rom[06066] = 16'h20a0;
  rom[06067] = 16'h30e1;
  rom[06068] = 16'h8b48;
  rom[06069] = 16'hedcd;
  rom[06070] = 16'hed89;
  rom[06071] = 16'hfdc9;
  rom[06072] = 16'hfd67;
  rom[06073] = 16'hfda8;
  rom[06074] = 16'hf587;
  rom[06075] = 16'hfda9;
  rom[06076] = 16'hfda8;
  rom[06077] = 16'hf5a9;
  rom[06078] = 16'hf5a8;
  rom[06079] = 16'hfda8;
  rom[06080] = 16'hfd88;
  rom[06081] = 16'hfda8;
  rom[06082] = 16'hf5a8;
  rom[06083] = 16'hfdc8;
  rom[06084] = 16'hfda8;
  rom[06085] = 16'hfdc8;
  rom[06086] = 16'hf5a9;
  rom[06087] = 16'hfdc9;
  rom[06088] = 16'hfda8;
  rom[06089] = 16'hfdc8;
  rom[06090] = 16'hf5a8;
  rom[06091] = 16'hfdc8;
  rom[06092] = 16'hfda8;
  rom[06093] = 16'hfdc9;
  rom[06094] = 16'hf5a9;
  rom[06095] = 16'hfdc9;
  rom[06096] = 16'hfda9;
  rom[06097] = 16'hfdc9;
  rom[06098] = 16'hf5a8;
  rom[06099] = 16'hfdc8;
  rom[06100] = 16'hfda8;
  rom[06101] = 16'hfdc8;
  rom[06102] = 16'hf5a9;
  rom[06103] = 16'hfdc8;
  rom[06104] = 16'hfda8;
  rom[06105] = 16'hfdc8;
  rom[06106] = 16'hf5a8;
  rom[06107] = 16'hfdc8;
  rom[06108] = 16'hfda8;
  rom[06109] = 16'hfdc8;
  rom[06110] = 16'hf5a8;
  rom[06111] = 16'hfdc8;
  rom[06112] = 16'hfd88;
  rom[06113] = 16'hfda9;
  rom[06114] = 16'hf589;
  rom[06115] = 16'hfda9;
  rom[06116] = 16'hfd89;
  rom[06117] = 16'hf5c8;
  rom[06118] = 16'hf5a7;
  rom[06119] = 16'hfda8;
  rom[06120] = 16'hfd88;
  rom[06121] = 16'hfd88;
  rom[06122] = 16'hf5a9;
  rom[06123] = 16'hf5ca;
  rom[06124] = 16'hd54b;
  rom[06125] = 16'h6244;
  rom[06126] = 16'h18a0;
  rom[06127] = 16'h18a1;
  rom[06128] = 16'h18a1;
  rom[06129] = 16'h18a2;
  rom[06130] = 16'h10a2;
  rom[06131] = 16'h10a3;
  rom[06132] = 16'h10a3;
  rom[06133] = 16'h18a3;
  rom[06134] = 16'h10c2;
  rom[06135] = 16'h18c3;
  rom[06136] = 16'h10a2;
  rom[06137] = 16'h10a2;
  rom[06138] = 16'h18e3;
  rom[06139] = 16'h94b2;
  rom[06140] = 16'hffdf;
  rom[06141] = 16'hffff;
  rom[06142] = 16'hffff;
  rom[06143] = 16'hffff;
  rom[06144] = 16'hffff;
  rom[06145] = 16'hffff;
  rom[06146] = 16'hffff;
  rom[06147] = 16'hffff;
  rom[06148] = 16'hffff;
  rom[06149] = 16'hffff;
  rom[06150] = 16'hffff;
  rom[06151] = 16'hffff;
  rom[06152] = 16'hffff;
  rom[06153] = 16'hffff;
  rom[06154] = 16'hffff;
  rom[06155] = 16'hffff;
  rom[06156] = 16'hffff;
  rom[06157] = 16'hffff;
  rom[06158] = 16'hffff;
  rom[06159] = 16'hffff;
  rom[06160] = 16'hffff;
  rom[06161] = 16'hffff;
  rom[06162] = 16'hffff;
  rom[06163] = 16'hffff;
  rom[06164] = 16'hffff;
  rom[06165] = 16'hffff;
  rom[06166] = 16'hffff;
  rom[06167] = 16'hffff;
  rom[06168] = 16'hffff;
  rom[06169] = 16'hffff;
  rom[06170] = 16'hffff;
  rom[06171] = 16'hffff;
  rom[06172] = 16'hffff;
  rom[06173] = 16'hffff;
  rom[06174] = 16'hffff;
  rom[06175] = 16'hffff;
  rom[06176] = 16'hffff;
  rom[06177] = 16'hffff;
  rom[06178] = 16'hffff;
  rom[06179] = 16'hffff;
  rom[06180] = 16'hffff;
  rom[06181] = 16'hffff;
  rom[06182] = 16'hffff;
  rom[06183] = 16'hffff;
  rom[06184] = 16'hffff;
  rom[06185] = 16'hffff;
  rom[06186] = 16'hffff;
  rom[06187] = 16'hffff;
  rom[06188] = 16'hffff;
  rom[06189] = 16'hffff;
  rom[06190] = 16'hffff;
  rom[06191] = 16'hffff;
  rom[06192] = 16'hffff;
  rom[06193] = 16'hffff;
  rom[06194] = 16'hffff;
  rom[06195] = 16'hffff;
  rom[06196] = 16'hffff;
  rom[06197] = 16'hffff;
  rom[06198] = 16'hffff;
  rom[06199] = 16'hffff;
  rom[06200] = 16'hffff;
  rom[06201] = 16'hffff;
  rom[06202] = 16'hffff;
  rom[06203] = 16'hffff;
  rom[06204] = 16'hffff;
  rom[06205] = 16'hffff;
  rom[06206] = 16'hffff;
  rom[06207] = 16'hffff;
  rom[06208] = 16'hffff;
  rom[06209] = 16'hffff;
  rom[06210] = 16'hffff;
  rom[06211] = 16'hffff;
  rom[06212] = 16'hffff;
  rom[06213] = 16'hffff;
  rom[06214] = 16'hffff;
  rom[06215] = 16'hffff;
  rom[06216] = 16'hffff;
  rom[06217] = 16'hffff;
  rom[06218] = 16'hffff;
  rom[06219] = 16'hffff;
  rom[06220] = 16'hffff;
  rom[06221] = 16'hffff;
  rom[06222] = 16'hffff;
  rom[06223] = 16'hffff;
  rom[06224] = 16'hffff;
  rom[06225] = 16'hffff;
  rom[06226] = 16'hffff;
  rom[06227] = 16'hffff;
  rom[06228] = 16'hffff;
  rom[06229] = 16'hffff;
  rom[06230] = 16'hffff;
  rom[06231] = 16'hffff;
  rom[06232] = 16'hffff;
  rom[06233] = 16'hffff;
  rom[06234] = 16'hffff;
  rom[06235] = 16'hffff;
  rom[06236] = 16'hffff;
  rom[06237] = 16'hffff;
  rom[06238] = 16'hffff;
  rom[06239] = 16'hffff;
  rom[06240] = 16'hffff;
  rom[06241] = 16'hffff;
  rom[06242] = 16'hffff;
  rom[06243] = 16'hffff;
  rom[06244] = 16'hffff;
  rom[06245] = 16'hffff;
  rom[06246] = 16'hffff;
  rom[06247] = 16'hffff;
  rom[06248] = 16'hffff;
  rom[06249] = 16'hffff;
  rom[06250] = 16'hffff;
  rom[06251] = 16'hffff;
  rom[06252] = 16'hffff;
  rom[06253] = 16'hffff;
  rom[06254] = 16'hef7d;
  rom[06255] = 16'h5aeb;
  rom[06256] = 16'h18e2;
  rom[06257] = 16'h18e2;
  rom[06258] = 16'h18c2;
  rom[06259] = 16'h18a2;
  rom[06260] = 16'h18a3;
  rom[06261] = 16'h18a3;
  rom[06262] = 16'h18a4;
  rom[06263] = 16'h1083;
  rom[06264] = 16'h1883;
  rom[06265] = 16'h18a2;
  rom[06266] = 16'h20e2;
  rom[06267] = 16'h2080;
  rom[06268] = 16'h82e7;
  rom[06269] = 16'he58c;
  rom[06270] = 16'hed89;
  rom[06271] = 16'hfd88;
  rom[06272] = 16'hfd87;
  rom[06273] = 16'hfda7;
  rom[06274] = 16'hfda8;
  rom[06275] = 16'hf5a9;
  rom[06276] = 16'hfdaa;
  rom[06277] = 16'hf5a9;
  rom[06278] = 16'hfda9;
  rom[06279] = 16'hfd88;
  rom[06280] = 16'hfda9;
  rom[06281] = 16'hfda8;
  rom[06282] = 16'hfdc9;
  rom[06283] = 16'hfda8;
  rom[06284] = 16'hfdc9;
  rom[06285] = 16'hfda8;
  rom[06286] = 16'hfdca;
  rom[06287] = 16'hfda9;
  rom[06288] = 16'hfdc9;
  rom[06289] = 16'hfda8;
  rom[06290] = 16'hfdc9;
  rom[06291] = 16'hfda8;
  rom[06292] = 16'hfdc9;
  rom[06293] = 16'hfda9;
  rom[06294] = 16'hfdca;
  rom[06295] = 16'hfda9;
  rom[06296] = 16'hfdca;
  rom[06297] = 16'hfda8;
  rom[06298] = 16'hfdc9;
  rom[06299] = 16'hfda8;
  rom[06300] = 16'hfde9;
  rom[06301] = 16'hfdc8;
  rom[06302] = 16'hfdc9;
  rom[06303] = 16'hfda8;
  rom[06304] = 16'hfdc9;
  rom[06305] = 16'hfda8;
  rom[06306] = 16'hfdc9;
  rom[06307] = 16'hfda8;
  rom[06308] = 16'hfdc9;
  rom[06309] = 16'hfda8;
  rom[06310] = 16'hfdc9;
  rom[06311] = 16'hfda8;
  rom[06312] = 16'hfdc9;
  rom[06313] = 16'hfda8;
  rom[06314] = 16'hfda9;
  rom[06315] = 16'hfd89;
  rom[06316] = 16'hfdaa;
  rom[06317] = 16'hf5a9;
  rom[06318] = 16'hfda8;
  rom[06319] = 16'hfd87;
  rom[06320] = 16'hfda8;
  rom[06321] = 16'hfd89;
  rom[06322] = 16'hfdca;
  rom[06323] = 16'hedaa;
  rom[06324] = 16'hd52c;
  rom[06325] = 16'h4982;
  rom[06326] = 16'h18c2;
  rom[06327] = 16'h18c2;
  rom[06328] = 16'h18c2;
  rom[06329] = 16'h18a2;
  rom[06330] = 16'h18a2;
  rom[06331] = 16'h10a2;
  rom[06332] = 16'h18a3;
  rom[06333] = 16'h18a3;
  rom[06334] = 16'h10c2;
  rom[06335] = 16'h10a2;
  rom[06336] = 16'h18c3;
  rom[06337] = 16'h10a2;
  rom[06338] = 16'h18e3;
  rom[06339] = 16'hc5f7;
  rom[06340] = 16'hffff;
  rom[06341] = 16'hffff;
  rom[06342] = 16'hffff;
  rom[06343] = 16'hffff;
  rom[06344] = 16'hffff;
  rom[06345] = 16'hffff;
  rom[06346] = 16'hffff;
  rom[06347] = 16'hffff;
  rom[06348] = 16'hffff;
  rom[06349] = 16'hffff;
  rom[06350] = 16'hffff;
  rom[06351] = 16'hffff;
  rom[06352] = 16'hffff;
  rom[06353] = 16'hffff;
  rom[06354] = 16'hffff;
  rom[06355] = 16'hffff;
  rom[06356] = 16'hffff;
  rom[06357] = 16'hffff;
  rom[06358] = 16'hffff;
  rom[06359] = 16'hffff;
  rom[06360] = 16'hffff;
  rom[06361] = 16'hffff;
  rom[06362] = 16'hffff;
  rom[06363] = 16'hffff;
  rom[06364] = 16'hffff;
  rom[06365] = 16'hffff;
  rom[06366] = 16'hffff;
  rom[06367] = 16'hffff;
  rom[06368] = 16'hffff;
  rom[06369] = 16'hffff;
  rom[06370] = 16'hffff;
  rom[06371] = 16'hffff;
  rom[06372] = 16'hffff;
  rom[06373] = 16'hffff;
  rom[06374] = 16'hffff;
  rom[06375] = 16'hffff;
  rom[06376] = 16'hffff;
  rom[06377] = 16'hffff;
  rom[06378] = 16'hffff;
  rom[06379] = 16'hffff;
  rom[06380] = 16'hffff;
  rom[06381] = 16'hffff;
  rom[06382] = 16'hffff;
  rom[06383] = 16'hffff;
  rom[06384] = 16'hffff;
  rom[06385] = 16'hffff;
  rom[06386] = 16'hffff;
  rom[06387] = 16'hffff;
  rom[06388] = 16'hffff;
  rom[06389] = 16'hffff;
  rom[06390] = 16'hffff;
  rom[06391] = 16'hffff;
  rom[06392] = 16'hffff;
  rom[06393] = 16'hffff;
  rom[06394] = 16'hffff;
  rom[06395] = 16'hffff;
  rom[06396] = 16'hffff;
  rom[06397] = 16'hffff;
  rom[06398] = 16'hffff;
  rom[06399] = 16'hffff;
  rom[06400] = 16'hffff;
  rom[06401] = 16'hffff;
  rom[06402] = 16'hffff;
  rom[06403] = 16'hffff;
  rom[06404] = 16'hffff;
  rom[06405] = 16'hffff;
  rom[06406] = 16'hffff;
  rom[06407] = 16'hffff;
  rom[06408] = 16'hffff;
  rom[06409] = 16'hffff;
  rom[06410] = 16'hffff;
  rom[06411] = 16'hffff;
  rom[06412] = 16'hffff;
  rom[06413] = 16'hffff;
  rom[06414] = 16'hffff;
  rom[06415] = 16'hffff;
  rom[06416] = 16'hffff;
  rom[06417] = 16'hffff;
  rom[06418] = 16'hffff;
  rom[06419] = 16'hffff;
  rom[06420] = 16'hffff;
  rom[06421] = 16'hffff;
  rom[06422] = 16'hffff;
  rom[06423] = 16'hffff;
  rom[06424] = 16'hffff;
  rom[06425] = 16'hffff;
  rom[06426] = 16'hffff;
  rom[06427] = 16'hffff;
  rom[06428] = 16'hffff;
  rom[06429] = 16'hffff;
  rom[06430] = 16'hffff;
  rom[06431] = 16'hffff;
  rom[06432] = 16'hffff;
  rom[06433] = 16'hffff;
  rom[06434] = 16'hffff;
  rom[06435] = 16'hffff;
  rom[06436] = 16'hffff;
  rom[06437] = 16'hffff;
  rom[06438] = 16'hffff;
  rom[06439] = 16'hffff;
  rom[06440] = 16'hffff;
  rom[06441] = 16'hffff;
  rom[06442] = 16'hffff;
  rom[06443] = 16'hffff;
  rom[06444] = 16'hffff;
  rom[06445] = 16'hffff;
  rom[06446] = 16'hffff;
  rom[06447] = 16'hffff;
  rom[06448] = 16'hffff;
  rom[06449] = 16'hffff;
  rom[06450] = 16'hffff;
  rom[06451] = 16'hffff;
  rom[06452] = 16'hffff;
  rom[06453] = 16'hffff;
  rom[06454] = 16'hffdf;
  rom[06455] = 16'h8c71;
  rom[06456] = 16'h18c2;
  rom[06457] = 16'h10a2;
  rom[06458] = 16'h10a2;
  rom[06459] = 16'h18c2;
  rom[06460] = 16'h10a1;
  rom[06461] = 16'h10a2;
  rom[06462] = 16'h10a2;
  rom[06463] = 16'h18c3;
  rom[06464] = 16'h0862;
  rom[06465] = 16'h18c3;
  rom[06466] = 16'h18c2;
  rom[06467] = 16'h20a1;
  rom[06468] = 16'h51c3;
  rom[06469] = 16'hd54c;
  rom[06470] = 16'hedaa;
  rom[06471] = 16'hfda9;
  rom[06472] = 16'hf587;
  rom[06473] = 16'hfdc8;
  rom[06474] = 16'hf587;
  rom[06475] = 16'hf589;
  rom[06476] = 16'hf5a9;
  rom[06477] = 16'hfda9;
  rom[06478] = 16'hfd88;
  rom[06479] = 16'hfdc8;
  rom[06480] = 16'hf5a8;
  rom[06481] = 16'hfdc8;
  rom[06482] = 16'hfda8;
  rom[06483] = 16'hfdc8;
  rom[06484] = 16'hf5a8;
  rom[06485] = 16'hfdc9;
  rom[06486] = 16'hfda9;
  rom[06487] = 16'hfdc9;
  rom[06488] = 16'hf5a8;
  rom[06489] = 16'hfdc8;
  rom[06490] = 16'hfda8;
  rom[06491] = 16'hfdc9;
  rom[06492] = 16'hf5c9;
  rom[06493] = 16'hfde9;
  rom[06494] = 16'hfdc9;
  rom[06495] = 16'hfde9;
  rom[06496] = 16'hf5c9;
  rom[06497] = 16'hfde9;
  rom[06498] = 16'hfdc9;
  rom[06499] = 16'hfde8;
  rom[06500] = 16'hf5c8;
  rom[06501] = 16'hfde8;
  rom[06502] = 16'hfdc9;
  rom[06503] = 16'hfde8;
  rom[06504] = 16'hf5a8;
  rom[06505] = 16'hfdc8;
  rom[06506] = 16'hfda8;
  rom[06507] = 16'hfdc8;
  rom[06508] = 16'hf5a8;
  rom[06509] = 16'hfdc8;
  rom[06510] = 16'hfda8;
  rom[06511] = 16'hfdc8;
  rom[06512] = 16'hf5a8;
  rom[06513] = 16'hfdc8;
  rom[06514] = 16'hfda9;
  rom[06515] = 16'hfdaa;
  rom[06516] = 16'hf589;
  rom[06517] = 16'hf5a9;
  rom[06518] = 16'hfda7;
  rom[06519] = 16'hfdc7;
  rom[06520] = 16'hfd87;
  rom[06521] = 16'hfd88;
  rom[06522] = 16'hed8a;
  rom[06523] = 16'he5cc;
  rom[06524] = 16'h9bc7;
  rom[06525] = 16'h3921;
  rom[06526] = 16'h10a2;
  rom[06527] = 16'h10c3;
  rom[06528] = 16'h10a2;
  rom[06529] = 16'h18c2;
  rom[06530] = 16'h10a2;
  rom[06531] = 16'h18a2;
  rom[06532] = 16'h18a3;
  rom[06533] = 16'h18a3;
  rom[06534] = 16'h10a2;
  rom[06535] = 16'h18a2;
  rom[06536] = 16'h10a2;
  rom[06537] = 16'h18a2;
  rom[06538] = 16'h4a28;
  rom[06539] = 16'he6fb;
  rom[06540] = 16'hffff;
  rom[06541] = 16'hffff;
  rom[06542] = 16'hffff;
  rom[06543] = 16'hffff;
  rom[06544] = 16'hffff;
  rom[06545] = 16'hffff;
  rom[06546] = 16'hffff;
  rom[06547] = 16'hffff;
  rom[06548] = 16'hffff;
  rom[06549] = 16'hffff;
  rom[06550] = 16'hffff;
  rom[06551] = 16'hffff;
  rom[06552] = 16'hffff;
  rom[06553] = 16'hffff;
  rom[06554] = 16'hffff;
  rom[06555] = 16'hffff;
  rom[06556] = 16'hffff;
  rom[06557] = 16'hffff;
  rom[06558] = 16'hffff;
  rom[06559] = 16'hffff;
  rom[06560] = 16'hffff;
  rom[06561] = 16'hffff;
  rom[06562] = 16'hffff;
  rom[06563] = 16'hffff;
  rom[06564] = 16'hffff;
  rom[06565] = 16'hffff;
  rom[06566] = 16'hffff;
  rom[06567] = 16'hffff;
  rom[06568] = 16'hffff;
  rom[06569] = 16'hffff;
  rom[06570] = 16'hffff;
  rom[06571] = 16'hffff;
  rom[06572] = 16'hffff;
  rom[06573] = 16'hffff;
  rom[06574] = 16'hffff;
  rom[06575] = 16'hffff;
  rom[06576] = 16'hffff;
  rom[06577] = 16'hffff;
  rom[06578] = 16'hffff;
  rom[06579] = 16'hffff;
  rom[06580] = 16'hffff;
  rom[06581] = 16'hffff;
  rom[06582] = 16'hffff;
  rom[06583] = 16'hffff;
  rom[06584] = 16'hffff;
  rom[06585] = 16'hffff;
  rom[06586] = 16'hffff;
  rom[06587] = 16'hffff;
  rom[06588] = 16'hffff;
  rom[06589] = 16'hffff;
  rom[06590] = 16'hffff;
  rom[06591] = 16'hffff;
  rom[06592] = 16'hffff;
  rom[06593] = 16'hffff;
  rom[06594] = 16'hffff;
  rom[06595] = 16'hffff;
  rom[06596] = 16'hffff;
  rom[06597] = 16'hffff;
  rom[06598] = 16'hffff;
  rom[06599] = 16'hffff;
  rom[06600] = 16'hffff;
  rom[06601] = 16'hffff;
  rom[06602] = 16'hffff;
  rom[06603] = 16'hffff;
  rom[06604] = 16'hffff;
  rom[06605] = 16'hffff;
  rom[06606] = 16'hffff;
  rom[06607] = 16'hffff;
  rom[06608] = 16'hffff;
  rom[06609] = 16'hffff;
  rom[06610] = 16'hffff;
  rom[06611] = 16'hffff;
  rom[06612] = 16'hffff;
  rom[06613] = 16'hffff;
  rom[06614] = 16'hffff;
  rom[06615] = 16'hffff;
  rom[06616] = 16'hffff;
  rom[06617] = 16'hffff;
  rom[06618] = 16'hffff;
  rom[06619] = 16'hffff;
  rom[06620] = 16'hffff;
  rom[06621] = 16'hffff;
  rom[06622] = 16'hffff;
  rom[06623] = 16'hffff;
  rom[06624] = 16'hffff;
  rom[06625] = 16'hffff;
  rom[06626] = 16'hffff;
  rom[06627] = 16'hffff;
  rom[06628] = 16'hffff;
  rom[06629] = 16'hffff;
  rom[06630] = 16'hffff;
  rom[06631] = 16'hffff;
  rom[06632] = 16'hffff;
  rom[06633] = 16'hffff;
  rom[06634] = 16'hffff;
  rom[06635] = 16'hffff;
  rom[06636] = 16'hffff;
  rom[06637] = 16'hffff;
  rom[06638] = 16'hffff;
  rom[06639] = 16'hffff;
  rom[06640] = 16'hffff;
  rom[06641] = 16'hffff;
  rom[06642] = 16'hffff;
  rom[06643] = 16'hffff;
  rom[06644] = 16'hffff;
  rom[06645] = 16'hffff;
  rom[06646] = 16'hffff;
  rom[06647] = 16'hffff;
  rom[06648] = 16'hffff;
  rom[06649] = 16'hffff;
  rom[06650] = 16'hffff;
  rom[06651] = 16'hffff;
  rom[06652] = 16'hffff;
  rom[06653] = 16'hffff;
  rom[06654] = 16'hffff;
  rom[06655] = 16'hc618;
  rom[06656] = 16'h3146;
  rom[06657] = 16'h10a3;
  rom[06658] = 16'h18a2;
  rom[06659] = 16'h18a2;
  rom[06660] = 16'h18c2;
  rom[06661] = 16'h10c2;
  rom[06662] = 16'h10c2;
  rom[06663] = 16'h10e2;
  rom[06664] = 16'h10a2;
  rom[06665] = 16'h10a2;
  rom[06666] = 16'h18c3;
  rom[06667] = 16'h18a2;
  rom[06668] = 16'h4122;
  rom[06669] = 16'hbcaa;
  rom[06670] = 16'hf5cd;
  rom[06671] = 16'hf56a;
  rom[06672] = 16'hfda9;
  rom[06673] = 16'hfd88;
  rom[06674] = 16'hfdca;
  rom[06675] = 16'hf589;
  rom[06676] = 16'hfdca;
  rom[06677] = 16'hfda9;
  rom[06678] = 16'hfdca;
  rom[06679] = 16'hfda8;
  rom[06680] = 16'hfdc9;
  rom[06681] = 16'hfda8;
  rom[06682] = 16'hfdc9;
  rom[06683] = 16'hfda8;
  rom[06684] = 16'hfdc9;
  rom[06685] = 16'hfda9;
  rom[06686] = 16'hfdca;
  rom[06687] = 16'hfda9;
  rom[06688] = 16'hfdc9;
  rom[06689] = 16'hfda8;
  rom[06690] = 16'hfde9;
  rom[06691] = 16'hfdc9;
  rom[06692] = 16'hfdea;
  rom[06693] = 16'hfdc9;
  rom[06694] = 16'hfdea;
  rom[06695] = 16'hfdc9;
  rom[06696] = 16'hfdea;
  rom[06697] = 16'hfdc9;
  rom[06698] = 16'hfdea;
  rom[06699] = 16'hfdc8;
  rom[06700] = 16'hfde9;
  rom[06701] = 16'hfdc8;
  rom[06702] = 16'hfdea;
  rom[06703] = 16'hfdc9;
  rom[06704] = 16'hfde9;
  rom[06705] = 16'hfda8;
  rom[06706] = 16'hfdea;
  rom[06707] = 16'hfda8;
  rom[06708] = 16'hfdc9;
  rom[06709] = 16'hfda8;
  rom[06710] = 16'hfdc9;
  rom[06711] = 16'hfda8;
  rom[06712] = 16'hfde9;
  rom[06713] = 16'hf5c7;
  rom[06714] = 16'hfdc9;
  rom[06715] = 16'hfda9;
  rom[06716] = 16'hfdaa;
  rom[06717] = 16'hf5a9;
  rom[06718] = 16'hfdc9;
  rom[06719] = 16'hfda7;
  rom[06720] = 16'hfd88;
  rom[06721] = 16'hfd89;
  rom[06722] = 16'hf5ab;
  rom[06723] = 16'hdd8d;
  rom[06724] = 16'h7ae5;
  rom[06725] = 16'h20c0;
  rom[06726] = 16'h18c3;
  rom[06727] = 16'h10c2;
  rom[06728] = 16'h18a2;
  rom[06729] = 16'h18a2;
  rom[06730] = 16'h18a3;
  rom[06731] = 16'h10a3;
  rom[06732] = 16'h18a3;
  rom[06733] = 16'h18a2;
  rom[06734] = 16'h18c2;
  rom[06735] = 16'h10a2;
  rom[06736] = 16'h18c2;
  rom[06737] = 16'h18c2;
  rom[06738] = 16'h7bae;
  rom[06739] = 16'hf77d;
  rom[06740] = 16'hffff;
  rom[06741] = 16'hffff;
  rom[06742] = 16'hffff;
  rom[06743] = 16'hffff;
  rom[06744] = 16'hffff;
  rom[06745] = 16'hffff;
  rom[06746] = 16'hffff;
  rom[06747] = 16'hffff;
  rom[06748] = 16'hffff;
  rom[06749] = 16'hffff;
  rom[06750] = 16'hffff;
  rom[06751] = 16'hffff;
  rom[06752] = 16'hffff;
  rom[06753] = 16'hffff;
  rom[06754] = 16'hffff;
  rom[06755] = 16'hffff;
  rom[06756] = 16'hffff;
  rom[06757] = 16'hffff;
  rom[06758] = 16'hffff;
  rom[06759] = 16'hffff;
  rom[06760] = 16'hffff;
  rom[06761] = 16'hffff;
  rom[06762] = 16'hffff;
  rom[06763] = 16'hffff;
  rom[06764] = 16'hffff;
  rom[06765] = 16'hffff;
  rom[06766] = 16'hffff;
  rom[06767] = 16'hffff;
  rom[06768] = 16'hffff;
  rom[06769] = 16'hffff;
  rom[06770] = 16'hffff;
  rom[06771] = 16'hffff;
  rom[06772] = 16'hffff;
  rom[06773] = 16'hffff;
  rom[06774] = 16'hffff;
  rom[06775] = 16'hffff;
  rom[06776] = 16'hffff;
  rom[06777] = 16'hffff;
  rom[06778] = 16'hffff;
  rom[06779] = 16'hffff;
  rom[06780] = 16'hffff;
  rom[06781] = 16'hffff;
  rom[06782] = 16'hffff;
  rom[06783] = 16'hffff;
  rom[06784] = 16'hffff;
  rom[06785] = 16'hffff;
  rom[06786] = 16'hffff;
  rom[06787] = 16'hffff;
  rom[06788] = 16'hffff;
  rom[06789] = 16'hffff;
  rom[06790] = 16'hffff;
  rom[06791] = 16'hffff;
  rom[06792] = 16'hffff;
  rom[06793] = 16'hffff;
  rom[06794] = 16'hffff;
  rom[06795] = 16'hffff;
  rom[06796] = 16'hffff;
  rom[06797] = 16'hffff;
  rom[06798] = 16'hffff;
  rom[06799] = 16'hffff;
  rom[06800] = 16'hffff;
  rom[06801] = 16'hffff;
  rom[06802] = 16'hffff;
  rom[06803] = 16'hffff;
  rom[06804] = 16'hffff;
  rom[06805] = 16'hffff;
  rom[06806] = 16'hffff;
  rom[06807] = 16'hffff;
  rom[06808] = 16'hffff;
  rom[06809] = 16'hffff;
  rom[06810] = 16'hffff;
  rom[06811] = 16'hffff;
  rom[06812] = 16'hffff;
  rom[06813] = 16'hffff;
  rom[06814] = 16'hffff;
  rom[06815] = 16'hffff;
  rom[06816] = 16'hffff;
  rom[06817] = 16'hffff;
  rom[06818] = 16'hffff;
  rom[06819] = 16'hffff;
  rom[06820] = 16'hffff;
  rom[06821] = 16'hffff;
  rom[06822] = 16'hffff;
  rom[06823] = 16'hffff;
  rom[06824] = 16'hffff;
  rom[06825] = 16'hffff;
  rom[06826] = 16'hffff;
  rom[06827] = 16'hffff;
  rom[06828] = 16'hffff;
  rom[06829] = 16'hffff;
  rom[06830] = 16'hffff;
  rom[06831] = 16'hffff;
  rom[06832] = 16'hffff;
  rom[06833] = 16'hffff;
  rom[06834] = 16'hffff;
  rom[06835] = 16'hffff;
  rom[06836] = 16'hffff;
  rom[06837] = 16'hffff;
  rom[06838] = 16'hffff;
  rom[06839] = 16'hffff;
  rom[06840] = 16'hffff;
  rom[06841] = 16'hffff;
  rom[06842] = 16'hffff;
  rom[06843] = 16'hffff;
  rom[06844] = 16'hffff;
  rom[06845] = 16'hffff;
  rom[06846] = 16'hffff;
  rom[06847] = 16'hffff;
  rom[06848] = 16'hffff;
  rom[06849] = 16'hffff;
  rom[06850] = 16'hffff;
  rom[06851] = 16'hffff;
  rom[06852] = 16'hffff;
  rom[06853] = 16'hffff;
  rom[06854] = 16'hffff;
  rom[06855] = 16'hef1c;
  rom[06856] = 16'h4a4a;
  rom[06857] = 16'h18a4;
  rom[06858] = 16'h1082;
  rom[06859] = 16'h18a3;
  rom[06860] = 16'h10a2;
  rom[06861] = 16'h18c3;
  rom[06862] = 16'h10c2;
  rom[06863] = 16'h10c3;
  rom[06864] = 16'h0882;
  rom[06865] = 16'h18e3;
  rom[06866] = 16'h10a2;
  rom[06867] = 16'h18c2;
  rom[06868] = 16'h20c1;
  rom[06869] = 16'h8347;
  rom[06870] = 16'hdd8c;
  rom[06871] = 16'hed8a;
  rom[06872] = 16'hfda9;
  rom[06873] = 16'hfd88;
  rom[06874] = 16'hf588;
  rom[06875] = 16'hfda8;
  rom[06876] = 16'hf588;
  rom[06877] = 16'hf5c9;
  rom[06878] = 16'hf5a9;
  rom[06879] = 16'hfdc8;
  rom[06880] = 16'hfda8;
  rom[06881] = 16'hfde8;
  rom[06882] = 16'hf5a8;
  rom[06883] = 16'hfdc8;
  rom[06884] = 16'hfda9;
  rom[06885] = 16'hfdc9;
  rom[06886] = 16'hf5a9;
  rom[06887] = 16'hfdc9;
  rom[06888] = 16'hfdc9;
  rom[06889] = 16'hfde9;
  rom[06890] = 16'hf5c9;
  rom[06891] = 16'hfde9;
  rom[06892] = 16'hfdc9;
  rom[06893] = 16'hfde9;
  rom[06894] = 16'hf5c9;
  rom[06895] = 16'hfde9;
  rom[06896] = 16'hfdc9;
  rom[06897] = 16'hfde9;
  rom[06898] = 16'hf5c9;
  rom[06899] = 16'hfde9;
  rom[06900] = 16'hfdc9;
  rom[06901] = 16'hfde9;
  rom[06902] = 16'hf5c9;
  rom[06903] = 16'hfde9;
  rom[06904] = 16'hfdc9;
  rom[06905] = 16'hfde9;
  rom[06906] = 16'hf5c9;
  rom[06907] = 16'hfde9;
  rom[06908] = 16'hfdc9;
  rom[06909] = 16'hfde9;
  rom[06910] = 16'hf5c8;
  rom[06911] = 16'hfde8;
  rom[06912] = 16'hf5c8;
  rom[06913] = 16'hf5e8;
  rom[06914] = 16'hf5a8;
  rom[06915] = 16'hfda8;
  rom[06916] = 16'hfd89;
  rom[06917] = 16'hfdc9;
  rom[06918] = 16'heda8;
  rom[06919] = 16'hfda8;
  rom[06920] = 16'hfda8;
  rom[06921] = 16'hfdaa;
  rom[06922] = 16'hed8b;
  rom[06923] = 16'hcd0c;
  rom[06924] = 16'h49a2;
  rom[06925] = 16'h20c1;
  rom[06926] = 16'h18a1;
  rom[06927] = 16'h18c2;
  rom[06928] = 16'h1082;
  rom[06929] = 16'h18a3;
  rom[06930] = 16'h1884;
  rom[06931] = 16'h18c4;
  rom[06932] = 16'h10a1;
  rom[06933] = 16'h10e2;
  rom[06934] = 16'h10a1;
  rom[06935] = 16'h18c2;
  rom[06936] = 16'h1081;
  rom[06937] = 16'h20e2;
  rom[06938] = 16'h5247;
  rom[06939] = 16'hc616;
  rom[06940] = 16'hffde;
  rom[06941] = 16'hffff;
  rom[06942] = 16'hffff;
  rom[06943] = 16'hffff;
  rom[06944] = 16'hffff;
  rom[06945] = 16'hffff;
  rom[06946] = 16'hffff;
  rom[06947] = 16'hffff;
  rom[06948] = 16'hffff;
  rom[06949] = 16'hffff;
  rom[06950] = 16'hffff;
  rom[06951] = 16'hffff;
  rom[06952] = 16'hffff;
  rom[06953] = 16'hffff;
  rom[06954] = 16'hffff;
  rom[06955] = 16'hffff;
  rom[06956] = 16'hffff;
  rom[06957] = 16'hffff;
  rom[06958] = 16'hffff;
  rom[06959] = 16'hffff;
  rom[06960] = 16'hffff;
  rom[06961] = 16'hffff;
  rom[06962] = 16'hffff;
  rom[06963] = 16'hffff;
  rom[06964] = 16'hffff;
  rom[06965] = 16'hffff;
  rom[06966] = 16'hffff;
  rom[06967] = 16'hffff;
  rom[06968] = 16'hffff;
  rom[06969] = 16'hffff;
  rom[06970] = 16'hffff;
  rom[06971] = 16'hffff;
  rom[06972] = 16'hffff;
  rom[06973] = 16'hffff;
  rom[06974] = 16'hffff;
  rom[06975] = 16'hffff;
  rom[06976] = 16'hffff;
  rom[06977] = 16'hffff;
  rom[06978] = 16'hffff;
  rom[06979] = 16'hffff;
  rom[06980] = 16'hffff;
  rom[06981] = 16'hffff;
  rom[06982] = 16'hffff;
  rom[06983] = 16'hffff;
  rom[06984] = 16'hffff;
  rom[06985] = 16'hffff;
  rom[06986] = 16'hffff;
  rom[06987] = 16'hffff;
  rom[06988] = 16'hffff;
  rom[06989] = 16'hffff;
  rom[06990] = 16'hffff;
  rom[06991] = 16'hffff;
  rom[06992] = 16'hffff;
  rom[06993] = 16'hffff;
  rom[06994] = 16'hffff;
  rom[06995] = 16'hffff;
  rom[06996] = 16'hffff;
  rom[06997] = 16'hffff;
  rom[06998] = 16'hffff;
  rom[06999] = 16'hffff;
  rom[07000] = 16'hffff;
  rom[07001] = 16'hffff;
  rom[07002] = 16'hffff;
  rom[07003] = 16'hffff;
  rom[07004] = 16'hffff;
  rom[07005] = 16'hffff;
  rom[07006] = 16'hffff;
  rom[07007] = 16'hffff;
  rom[07008] = 16'hffff;
  rom[07009] = 16'hffff;
  rom[07010] = 16'hffff;
  rom[07011] = 16'hffff;
  rom[07012] = 16'hffff;
  rom[07013] = 16'hffff;
  rom[07014] = 16'hffff;
  rom[07015] = 16'hffff;
  rom[07016] = 16'hffff;
  rom[07017] = 16'hffff;
  rom[07018] = 16'hffff;
  rom[07019] = 16'hffff;
  rom[07020] = 16'hffff;
  rom[07021] = 16'hffff;
  rom[07022] = 16'hffff;
  rom[07023] = 16'hffff;
  rom[07024] = 16'hffff;
  rom[07025] = 16'hffff;
  rom[07026] = 16'hffff;
  rom[07027] = 16'hffff;
  rom[07028] = 16'hffff;
  rom[07029] = 16'hffff;
  rom[07030] = 16'hffff;
  rom[07031] = 16'hffff;
  rom[07032] = 16'hffff;
  rom[07033] = 16'hffff;
  rom[07034] = 16'hffff;
  rom[07035] = 16'hffff;
  rom[07036] = 16'hffff;
  rom[07037] = 16'hffff;
  rom[07038] = 16'hffff;
  rom[07039] = 16'hffff;
  rom[07040] = 16'hffff;
  rom[07041] = 16'hffff;
  rom[07042] = 16'hffff;
  rom[07043] = 16'hffff;
  rom[07044] = 16'hffff;
  rom[07045] = 16'hffff;
  rom[07046] = 16'hffff;
  rom[07047] = 16'hffff;
  rom[07048] = 16'hffff;
  rom[07049] = 16'hffff;
  rom[07050] = 16'hffff;
  rom[07051] = 16'hffff;
  rom[07052] = 16'hffff;
  rom[07053] = 16'hffff;
  rom[07054] = 16'hffff;
  rom[07055] = 16'hf77e;
  rom[07056] = 16'h83d0;
  rom[07057] = 16'h28e4;
  rom[07058] = 16'h18a3;
  rom[07059] = 16'h10a2;
  rom[07060] = 16'h18c3;
  rom[07061] = 16'h10a2;
  rom[07062] = 16'h10c3;
  rom[07063] = 16'h10c2;
  rom[07064] = 16'h10a2;
  rom[07065] = 16'h18c2;
  rom[07066] = 16'h18a2;
  rom[07067] = 16'h18a2;
  rom[07068] = 16'h20a1;
  rom[07069] = 16'h5203;
  rom[07070] = 16'hcd2d;
  rom[07071] = 16'he5ab;
  rom[07072] = 16'hfdaa;
  rom[07073] = 16'hfda8;
  rom[07074] = 16'hfda9;
  rom[07075] = 16'hfda8;
  rom[07076] = 16'hfdc9;
  rom[07077] = 16'hf5ca;
  rom[07078] = 16'hf5ca;
  rom[07079] = 16'hfdc8;
  rom[07080] = 16'hfde9;
  rom[07081] = 16'hfdc8;
  rom[07082] = 16'hfde9;
  rom[07083] = 16'hfdc8;
  rom[07084] = 16'hfdea;
  rom[07085] = 16'hfdc9;
  rom[07086] = 16'hfdea;
  rom[07087] = 16'hfdc9;
  rom[07088] = 16'hfde9;
  rom[07089] = 16'hfdc9;
  rom[07090] = 16'hfdea;
  rom[07091] = 16'hfdc9;
  rom[07092] = 16'hfdea;
  rom[07093] = 16'hfdc9;
  rom[07094] = 16'hfdea;
  rom[07095] = 16'hfdc9;
  rom[07096] = 16'hfdea;
  rom[07097] = 16'hfdc9;
  rom[07098] = 16'hfdea;
  rom[07099] = 16'hfdc9;
  rom[07100] = 16'hfdea;
  rom[07101] = 16'hfdc9;
  rom[07102] = 16'hfdea;
  rom[07103] = 16'hfdc9;
  rom[07104] = 16'hfdea;
  rom[07105] = 16'hfdc9;
  rom[07106] = 16'hfdea;
  rom[07107] = 16'hfdc9;
  rom[07108] = 16'hfdea;
  rom[07109] = 16'hfdc9;
  rom[07110] = 16'hfde9;
  rom[07111] = 16'hfdc8;
  rom[07112] = 16'hf5e9;
  rom[07113] = 16'hf5c9;
  rom[07114] = 16'hfdc9;
  rom[07115] = 16'hfda8;
  rom[07116] = 16'hfda9;
  rom[07117] = 16'hf5a9;
  rom[07118] = 16'hf5c9;
  rom[07119] = 16'hfdc8;
  rom[07120] = 16'hfd89;
  rom[07121] = 16'hfd8a;
  rom[07122] = 16'hed8c;
  rom[07123] = 16'ha429;
  rom[07124] = 16'h28c1;
  rom[07125] = 16'h20a1;
  rom[07126] = 16'h18a2;
  rom[07127] = 16'h10a2;
  rom[07128] = 16'h18c3;
  rom[07129] = 16'h20a3;
  rom[07130] = 16'h18a4;
  rom[07131] = 16'h10a3;
  rom[07132] = 16'h10e2;
  rom[07133] = 16'h10c1;
  rom[07134] = 16'h18c2;
  rom[07135] = 16'h18a2;
  rom[07136] = 16'h20c3;
  rom[07137] = 16'h41a4;
  rom[07138] = 16'h9c2d;
  rom[07139] = 16'h7349;
  rom[07140] = 16'hd677;
  rom[07141] = 16'hffdf;
  rom[07142] = 16'hffff;
  rom[07143] = 16'hffdf;
  rom[07144] = 16'hffff;
  rom[07145] = 16'hffff;
  rom[07146] = 16'hffff;
  rom[07147] = 16'hffff;
  rom[07148] = 16'hffff;
  rom[07149] = 16'hffff;
  rom[07150] = 16'hffff;
  rom[07151] = 16'hffff;
  rom[07152] = 16'hffff;
  rom[07153] = 16'hffff;
  rom[07154] = 16'hffff;
  rom[07155] = 16'hffff;
  rom[07156] = 16'hffff;
  rom[07157] = 16'hffff;
  rom[07158] = 16'hffff;
  rom[07159] = 16'hffff;
  rom[07160] = 16'hffff;
  rom[07161] = 16'hffff;
  rom[07162] = 16'hffff;
  rom[07163] = 16'hffff;
  rom[07164] = 16'hffff;
  rom[07165] = 16'hffff;
  rom[07166] = 16'hffff;
  rom[07167] = 16'hffff;
  rom[07168] = 16'hffff;
  rom[07169] = 16'hffff;
  rom[07170] = 16'hffff;
  rom[07171] = 16'hffff;
  rom[07172] = 16'hffff;
  rom[07173] = 16'hffff;
  rom[07174] = 16'hffff;
  rom[07175] = 16'hffff;
  rom[07176] = 16'hffff;
  rom[07177] = 16'hffff;
  rom[07178] = 16'hffff;
  rom[07179] = 16'hffff;
  rom[07180] = 16'hffff;
  rom[07181] = 16'hffff;
  rom[07182] = 16'hffff;
  rom[07183] = 16'hffff;
  rom[07184] = 16'hffff;
  rom[07185] = 16'hffff;
  rom[07186] = 16'hffff;
  rom[07187] = 16'hffff;
  rom[07188] = 16'hffff;
  rom[07189] = 16'hffff;
  rom[07190] = 16'hffff;
  rom[07191] = 16'hffff;
  rom[07192] = 16'hffff;
  rom[07193] = 16'hffff;
  rom[07194] = 16'hffff;
  rom[07195] = 16'hffff;
  rom[07196] = 16'hffff;
  rom[07197] = 16'hffff;
  rom[07198] = 16'hffff;
  rom[07199] = 16'hffff;
  rom[07200] = 16'hffff;
  rom[07201] = 16'hffff;
  rom[07202] = 16'hffff;
  rom[07203] = 16'hffff;
  rom[07204] = 16'hffff;
  rom[07205] = 16'hffff;
  rom[07206] = 16'hffff;
  rom[07207] = 16'hffff;
  rom[07208] = 16'hffff;
  rom[07209] = 16'hffff;
  rom[07210] = 16'hffff;
  rom[07211] = 16'hffff;
  rom[07212] = 16'hffff;
  rom[07213] = 16'hffff;
  rom[07214] = 16'hffff;
  rom[07215] = 16'hffff;
  rom[07216] = 16'hffff;
  rom[07217] = 16'hffff;
  rom[07218] = 16'hffff;
  rom[07219] = 16'hffff;
  rom[07220] = 16'hffff;
  rom[07221] = 16'hffff;
  rom[07222] = 16'hffff;
  rom[07223] = 16'hffff;
  rom[07224] = 16'hffff;
  rom[07225] = 16'hffff;
  rom[07226] = 16'hffff;
  rom[07227] = 16'hffff;
  rom[07228] = 16'hffff;
  rom[07229] = 16'hffff;
  rom[07230] = 16'hffff;
  rom[07231] = 16'hffff;
  rom[07232] = 16'hffff;
  rom[07233] = 16'hffff;
  rom[07234] = 16'hffff;
  rom[07235] = 16'hffff;
  rom[07236] = 16'hffff;
  rom[07237] = 16'hffff;
  rom[07238] = 16'hffff;
  rom[07239] = 16'hffff;
  rom[07240] = 16'hffff;
  rom[07241] = 16'hffff;
  rom[07242] = 16'hffff;
  rom[07243] = 16'hffff;
  rom[07244] = 16'hffff;
  rom[07245] = 16'hffff;
  rom[07246] = 16'hffff;
  rom[07247] = 16'hffff;
  rom[07248] = 16'hffff;
  rom[07249] = 16'hffff;
  rom[07250] = 16'hffff;
  rom[07251] = 16'hffff;
  rom[07252] = 16'hffff;
  rom[07253] = 16'hffbf;
  rom[07254] = 16'hffdf;
  rom[07255] = 16'hffdf;
  rom[07256] = 16'ha4d2;
  rom[07257] = 16'h1861;
  rom[07258] = 16'h1061;
  rom[07259] = 16'h18a3;
  rom[07260] = 16'h18c3;
  rom[07261] = 16'h18e4;
  rom[07262] = 16'h10c2;
  rom[07263] = 16'h18c2;
  rom[07264] = 16'h10a1;
  rom[07265] = 16'h18c2;
  rom[07266] = 16'h18a2;
  rom[07267] = 16'h18a2;
  rom[07268] = 16'h18a1;
  rom[07269] = 16'h3120;
  rom[07270] = 16'ha44a;
  rom[07271] = 16'hedcd;
  rom[07272] = 16'hf58a;
  rom[07273] = 16'hfdc9;
  rom[07274] = 16'hfd87;
  rom[07275] = 16'hfda8;
  rom[07276] = 16'hf588;
  rom[07277] = 16'hf5ca;
  rom[07278] = 16'hf5a9;
  rom[07279] = 16'hfdc8;
  rom[07280] = 16'hf5c8;
  rom[07281] = 16'hfde8;
  rom[07282] = 16'hfdc8;
  rom[07283] = 16'hfde8;
  rom[07284] = 16'hf5c8;
  rom[07285] = 16'hfde8;
  rom[07286] = 16'hfdc9;
  rom[07287] = 16'hfde8;
  rom[07288] = 16'hf5c8;
  rom[07289] = 16'hfde8;
  rom[07290] = 16'hfdc9;
  rom[07291] = 16'hfde9;
  rom[07292] = 16'hf5c9;
  rom[07293] = 16'hfde9;
  rom[07294] = 16'hfdc9;
  rom[07295] = 16'hfde9;
  rom[07296] = 16'hf5c9;
  rom[07297] = 16'hfde9;
  rom[07298] = 16'hfdc9;
  rom[07299] = 16'hfde9;
  rom[07300] = 16'hf5c9;
  rom[07301] = 16'hfde9;
  rom[07302] = 16'hfdc9;
  rom[07303] = 16'hfde9;
  rom[07304] = 16'hf5c9;
  rom[07305] = 16'hfde9;
  rom[07306] = 16'hfdc9;
  rom[07307] = 16'hfde9;
  rom[07308] = 16'hf5c9;
  rom[07309] = 16'hfde9;
  rom[07310] = 16'hfdc9;
  rom[07311] = 16'hfde9;
  rom[07312] = 16'hf5c9;
  rom[07313] = 16'hf5e9;
  rom[07314] = 16'hf5a9;
  rom[07315] = 16'hfdc8;
  rom[07316] = 16'hf5a8;
  rom[07317] = 16'hf5c8;
  rom[07318] = 16'hf5a8;
  rom[07319] = 16'hf588;
  rom[07320] = 16'hfd89;
  rom[07321] = 16'hfd8b;
  rom[07322] = 16'hdd2b;
  rom[07323] = 16'h8305;
  rom[07324] = 16'h18a0;
  rom[07325] = 16'h18a2;
  rom[07326] = 16'h18a2;
  rom[07327] = 16'h18c3;
  rom[07328] = 16'h1882;
  rom[07329] = 16'h18a3;
  rom[07330] = 16'h1883;
  rom[07331] = 16'h1082;
  rom[07332] = 16'h10a1;
  rom[07333] = 16'h10e1;
  rom[07334] = 16'h10a2;
  rom[07335] = 16'h18a3;
  rom[07336] = 16'h1881;
  rom[07337] = 16'h7b07;
  rom[07338] = 16'hd590;
  rom[07339] = 16'ha42b;
  rom[07340] = 16'h7309;
  rom[07341] = 16'heed9;
  rom[07342] = 16'hffde;
  rom[07343] = 16'hffff;
  rom[07344] = 16'hf7de;
  rom[07345] = 16'hffff;
  rom[07346] = 16'hffff;
  rom[07347] = 16'hffff;
  rom[07348] = 16'hffff;
  rom[07349] = 16'hffff;
  rom[07350] = 16'hffff;
  rom[07351] = 16'hffff;
  rom[07352] = 16'hffff;
  rom[07353] = 16'hffff;
  rom[07354] = 16'hffff;
  rom[07355] = 16'hffff;
  rom[07356] = 16'hffff;
  rom[07357] = 16'hffff;
  rom[07358] = 16'hffff;
  rom[07359] = 16'hffff;
  rom[07360] = 16'hffff;
  rom[07361] = 16'hffff;
  rom[07362] = 16'hffff;
  rom[07363] = 16'hffff;
  rom[07364] = 16'hffff;
  rom[07365] = 16'hffff;
  rom[07366] = 16'hffff;
  rom[07367] = 16'hffff;
  rom[07368] = 16'hffff;
  rom[07369] = 16'hffff;
  rom[07370] = 16'hffff;
  rom[07371] = 16'hffff;
  rom[07372] = 16'hffff;
  rom[07373] = 16'hffff;
  rom[07374] = 16'hffff;
  rom[07375] = 16'hffff;
  rom[07376] = 16'hffff;
  rom[07377] = 16'hffff;
  rom[07378] = 16'hffff;
  rom[07379] = 16'hffff;
  rom[07380] = 16'hffff;
  rom[07381] = 16'hffff;
  rom[07382] = 16'hffff;
  rom[07383] = 16'hffff;
  rom[07384] = 16'hffff;
  rom[07385] = 16'hffff;
  rom[07386] = 16'hffff;
  rom[07387] = 16'hffff;
  rom[07388] = 16'hffff;
  rom[07389] = 16'hffff;
  rom[07390] = 16'hffff;
  rom[07391] = 16'hffff;
  rom[07392] = 16'hffff;
  rom[07393] = 16'hffff;
  rom[07394] = 16'hffff;
  rom[07395] = 16'hffff;
  rom[07396] = 16'hffff;
  rom[07397] = 16'hffff;
  rom[07398] = 16'hffff;
  rom[07399] = 16'hffff;
  rom[07400] = 16'hffff;
  rom[07401] = 16'hffff;
  rom[07402] = 16'hffff;
  rom[07403] = 16'hffff;
  rom[07404] = 16'hffff;
  rom[07405] = 16'hffff;
  rom[07406] = 16'hffff;
  rom[07407] = 16'hffff;
  rom[07408] = 16'hffff;
  rom[07409] = 16'hffff;
  rom[07410] = 16'hffff;
  rom[07411] = 16'hffff;
  rom[07412] = 16'hffff;
  rom[07413] = 16'hffff;
  rom[07414] = 16'hffff;
  rom[07415] = 16'hffff;
  rom[07416] = 16'hffff;
  rom[07417] = 16'hffff;
  rom[07418] = 16'hffff;
  rom[07419] = 16'hffff;
  rom[07420] = 16'hffff;
  rom[07421] = 16'hffff;
  rom[07422] = 16'hffff;
  rom[07423] = 16'hffff;
  rom[07424] = 16'hffff;
  rom[07425] = 16'hffff;
  rom[07426] = 16'hffff;
  rom[07427] = 16'hffff;
  rom[07428] = 16'hffff;
  rom[07429] = 16'hffff;
  rom[07430] = 16'hffff;
  rom[07431] = 16'hffff;
  rom[07432] = 16'hffff;
  rom[07433] = 16'hffff;
  rom[07434] = 16'hffff;
  rom[07435] = 16'hffff;
  rom[07436] = 16'hffff;
  rom[07437] = 16'hffff;
  rom[07438] = 16'hffff;
  rom[07439] = 16'hffff;
  rom[07440] = 16'hffff;
  rom[07441] = 16'hffff;
  rom[07442] = 16'hffff;
  rom[07443] = 16'hffff;
  rom[07444] = 16'hffff;
  rom[07445] = 16'hffff;
  rom[07446] = 16'hffff;
  rom[07447] = 16'hffff;
  rom[07448] = 16'hffff;
  rom[07449] = 16'hffff;
  rom[07450] = 16'hffff;
  rom[07451] = 16'hffff;
  rom[07452] = 16'hffff;
  rom[07453] = 16'hffbf;
  rom[07454] = 16'hffbf;
  rom[07455] = 16'hbd95;
  rom[07456] = 16'h730a;
  rom[07457] = 16'h4183;
  rom[07458] = 16'h28c1;
  rom[07459] = 16'h20a2;
  rom[07460] = 16'h18a3;
  rom[07461] = 16'h10a3;
  rom[07462] = 16'h10a3;
  rom[07463] = 16'h10c2;
  rom[07464] = 16'h10a2;
  rom[07465] = 16'h18c2;
  rom[07466] = 16'h18a2;
  rom[07467] = 16'h18a2;
  rom[07468] = 16'h18c2;
  rom[07469] = 16'h1860;
  rom[07470] = 16'h7ae6;
  rom[07471] = 16'hdd8d;
  rom[07472] = 16'hf5cb;
  rom[07473] = 16'hf5c8;
  rom[07474] = 16'hfda8;
  rom[07475] = 16'hfda8;
  rom[07476] = 16'hfdc9;
  rom[07477] = 16'hf5c9;
  rom[07478] = 16'hf5ea;
  rom[07479] = 16'hfdc8;
  rom[07480] = 16'hfde9;
  rom[07481] = 16'hfdc8;
  rom[07482] = 16'hfde9;
  rom[07483] = 16'hfdc8;
  rom[07484] = 16'hfde9;
  rom[07485] = 16'hfde8;
  rom[07486] = 16'hfde9;
  rom[07487] = 16'hfde8;
  rom[07488] = 16'hfde9;
  rom[07489] = 16'hfdc8;
  rom[07490] = 16'hfde9;
  rom[07491] = 16'hfdc9;
  rom[07492] = 16'hfdea;
  rom[07493] = 16'hfdc9;
  rom[07494] = 16'hfdea;
  rom[07495] = 16'hfdc9;
  rom[07496] = 16'hfdea;
  rom[07497] = 16'hfdc9;
  rom[07498] = 16'hfdea;
  rom[07499] = 16'hfdc9;
  rom[07500] = 16'hfdea;
  rom[07501] = 16'hfdc9;
  rom[07502] = 16'hfdea;
  rom[07503] = 16'hfdc9;
  rom[07504] = 16'hfdea;
  rom[07505] = 16'hfdc9;
  rom[07506] = 16'hfdea;
  rom[07507] = 16'hfdc9;
  rom[07508] = 16'hfdea;
  rom[07509] = 16'hfdc9;
  rom[07510] = 16'hfdea;
  rom[07511] = 16'hfdc9;
  rom[07512] = 16'hfdea;
  rom[07513] = 16'hf5ca;
  rom[07514] = 16'hfdca;
  rom[07515] = 16'hfda9;
  rom[07516] = 16'hfdc9;
  rom[07517] = 16'hf5c8;
  rom[07518] = 16'hfde9;
  rom[07519] = 16'hf588;
  rom[07520] = 16'hfdaa;
  rom[07521] = 16'hf5ac;
  rom[07522] = 16'hccec;
  rom[07523] = 16'h49e2;
  rom[07524] = 16'h1881;
  rom[07525] = 16'h18a2;
  rom[07526] = 16'h18a3;
  rom[07527] = 16'h18a2;
  rom[07528] = 16'h18c2;
  rom[07529] = 16'h1882;
  rom[07530] = 16'h18a3;
  rom[07531] = 16'h1062;
  rom[07532] = 16'h18c3;
  rom[07533] = 16'h08a1;
  rom[07534] = 16'h20c3;
  rom[07535] = 16'h20a3;
  rom[07536] = 16'h3902;
  rom[07537] = 16'ha429;
  rom[07538] = 16'he58d;
  rom[07539] = 16'hdd2d;
  rom[07540] = 16'h9b89;
  rom[07541] = 16'h93ec;
  rom[07542] = 16'hf73b;
  rom[07543] = 16'hffde;
  rom[07544] = 16'hffdf;
  rom[07545] = 16'hffff;
  rom[07546] = 16'hffff;
  rom[07547] = 16'hffff;
  rom[07548] = 16'hffff;
  rom[07549] = 16'hffff;
  rom[07550] = 16'hffff;
  rom[07551] = 16'hffff;
  rom[07552] = 16'hffff;
  rom[07553] = 16'hffff;
  rom[07554] = 16'hffff;
  rom[07555] = 16'hffff;
  rom[07556] = 16'hffff;
  rom[07557] = 16'hffff;
  rom[07558] = 16'hffff;
  rom[07559] = 16'hffff;
  rom[07560] = 16'hffff;
  rom[07561] = 16'hffff;
  rom[07562] = 16'hffff;
  rom[07563] = 16'hffff;
  rom[07564] = 16'hffff;
  rom[07565] = 16'hffff;
  rom[07566] = 16'hffff;
  rom[07567] = 16'hffff;
  rom[07568] = 16'hffff;
  rom[07569] = 16'hffff;
  rom[07570] = 16'hffff;
  rom[07571] = 16'hffff;
  rom[07572] = 16'hffff;
  rom[07573] = 16'hffff;
  rom[07574] = 16'hffff;
  rom[07575] = 16'hffff;
  rom[07576] = 16'hffff;
  rom[07577] = 16'hffff;
  rom[07578] = 16'hffff;
  rom[07579] = 16'hffff;
  rom[07580] = 16'hffff;
  rom[07581] = 16'hffff;
  rom[07582] = 16'hffff;
  rom[07583] = 16'hffff;
  rom[07584] = 16'hffff;
  rom[07585] = 16'hffff;
  rom[07586] = 16'hffff;
  rom[07587] = 16'hffff;
  rom[07588] = 16'hffff;
  rom[07589] = 16'hffff;
  rom[07590] = 16'hffff;
  rom[07591] = 16'hffff;
  rom[07592] = 16'hffff;
  rom[07593] = 16'hffff;
  rom[07594] = 16'hffff;
  rom[07595] = 16'hffff;
  rom[07596] = 16'hffff;
  rom[07597] = 16'hffff;
  rom[07598] = 16'hffff;
  rom[07599] = 16'hffff;
  rom[07600] = 16'hffff;
  rom[07601] = 16'hffff;
  rom[07602] = 16'hffff;
  rom[07603] = 16'hffff;
  rom[07604] = 16'hffff;
  rom[07605] = 16'hffff;
  rom[07606] = 16'hffff;
  rom[07607] = 16'hffff;
  rom[07608] = 16'hffff;
  rom[07609] = 16'hffff;
  rom[07610] = 16'hffff;
  rom[07611] = 16'hffff;
  rom[07612] = 16'hffff;
  rom[07613] = 16'hffff;
  rom[07614] = 16'hffff;
  rom[07615] = 16'hffff;
  rom[07616] = 16'hffff;
  rom[07617] = 16'hffff;
  rom[07618] = 16'hffff;
  rom[07619] = 16'hffff;
  rom[07620] = 16'hffff;
  rom[07621] = 16'hffff;
  rom[07622] = 16'hffff;
  rom[07623] = 16'hffff;
  rom[07624] = 16'hffff;
  rom[07625] = 16'hffff;
  rom[07626] = 16'hffff;
  rom[07627] = 16'hffff;
  rom[07628] = 16'hffff;
  rom[07629] = 16'hffff;
  rom[07630] = 16'hffff;
  rom[07631] = 16'hffff;
  rom[07632] = 16'hffff;
  rom[07633] = 16'hffff;
  rom[07634] = 16'hffff;
  rom[07635] = 16'hffff;
  rom[07636] = 16'hffff;
  rom[07637] = 16'hffff;
  rom[07638] = 16'hffff;
  rom[07639] = 16'hffff;
  rom[07640] = 16'hffff;
  rom[07641] = 16'hffff;
  rom[07642] = 16'hffff;
  rom[07643] = 16'hffff;
  rom[07644] = 16'hffff;
  rom[07645] = 16'hffff;
  rom[07646] = 16'hffff;
  rom[07647] = 16'hffff;
  rom[07648] = 16'hffff;
  rom[07649] = 16'hffff;
  rom[07650] = 16'hffdf;
  rom[07651] = 16'hffff;
  rom[07652] = 16'hffdf;
  rom[07653] = 16'hffbe;
  rom[07654] = 16'hc5b4;
  rom[07655] = 16'h5a66;
  rom[07656] = 16'ha44c;
  rom[07657] = 16'h8349;
  rom[07658] = 16'h2880;
  rom[07659] = 16'h1882;
  rom[07660] = 16'h20c4;
  rom[07661] = 16'h1063;
  rom[07662] = 16'h10a3;
  rom[07663] = 16'h18c3;
  rom[07664] = 16'h18c2;
  rom[07665] = 16'h18c2;
  rom[07666] = 16'h1882;
  rom[07667] = 16'h18a3;
  rom[07668] = 16'h10a2;
  rom[07669] = 16'h20c1;
  rom[07670] = 16'h41a2;
  rom[07671] = 16'hc4ec;
  rom[07672] = 16'hedcb;
  rom[07673] = 16'hf5c8;
  rom[07674] = 16'hfda8;
  rom[07675] = 16'hfdc8;
  rom[07676] = 16'hfd89;
  rom[07677] = 16'hf5c9;
  rom[07678] = 16'heda8;
  rom[07679] = 16'hfde8;
  rom[07680] = 16'hfdc8;
  rom[07681] = 16'hfde8;
  rom[07682] = 16'hf5c8;
  rom[07683] = 16'hfde8;
  rom[07684] = 16'hfde8;
  rom[07685] = 16'hfe09;
  rom[07686] = 16'hf5e9;
  rom[07687] = 16'hfe09;
  rom[07688] = 16'hfde8;
  rom[07689] = 16'hfe08;
  rom[07690] = 16'hf5e9;
  rom[07691] = 16'hfe09;
  rom[07692] = 16'hfde9;
  rom[07693] = 16'hfe09;
  rom[07694] = 16'hf5e9;
  rom[07695] = 16'hfe09;
  rom[07696] = 16'hfde9;
  rom[07697] = 16'hfe09;
  rom[07698] = 16'hf5e9;
  rom[07699] = 16'hfe09;
  rom[07700] = 16'hfde9;
  rom[07701] = 16'hfe09;
  rom[07702] = 16'hf5e9;
  rom[07703] = 16'hfe09;
  rom[07704] = 16'hfde9;
  rom[07705] = 16'hfe09;
  rom[07706] = 16'hf5c9;
  rom[07707] = 16'hfde9;
  rom[07708] = 16'hfdc9;
  rom[07709] = 16'hfde9;
  rom[07710] = 16'hf5c9;
  rom[07711] = 16'hfde8;
  rom[07712] = 16'hfdc9;
  rom[07713] = 16'hfde9;
  rom[07714] = 16'hf5a9;
  rom[07715] = 16'hfdc9;
  rom[07716] = 16'hfdc8;
  rom[07717] = 16'hf5e8;
  rom[07718] = 16'hf5c7;
  rom[07719] = 16'hfdc8;
  rom[07720] = 16'hf569;
  rom[07721] = 16'hf58d;
  rom[07722] = 16'h93a8;
  rom[07723] = 16'h2901;
  rom[07724] = 16'h10a1;
  rom[07725] = 16'h18e4;
  rom[07726] = 16'h10e3;
  rom[07727] = 16'h10a2;
  rom[07728] = 16'h18c2;
  rom[07729] = 16'h1881;
  rom[07730] = 16'h1882;
  rom[07731] = 16'h1083;
  rom[07732] = 16'h10e3;
  rom[07733] = 16'h1082;
  rom[07734] = 16'h18c2;
  rom[07735] = 16'h1860;
  rom[07736] = 16'h5a24;
  rom[07737] = 16'hd54b;
  rom[07738] = 16'hed8a;
  rom[07739] = 16'hed6c;
  rom[07740] = 16'hccab;
  rom[07741] = 16'h9368;
  rom[07742] = 16'haccf;
  rom[07743] = 16'hfffe;
  rom[07744] = 16'hffbf;
  rom[07745] = 16'hffff;
  rom[07746] = 16'hffff;
  rom[07747] = 16'hffff;
  rom[07748] = 16'hffff;
  rom[07749] = 16'hffff;
  rom[07750] = 16'hffff;
  rom[07751] = 16'hffff;
  rom[07752] = 16'hffff;
  rom[07753] = 16'hffff;
  rom[07754] = 16'hffff;
  rom[07755] = 16'hffff;
  rom[07756] = 16'hffff;
  rom[07757] = 16'hffff;
  rom[07758] = 16'hffff;
  rom[07759] = 16'hffff;
  rom[07760] = 16'hffff;
  rom[07761] = 16'hffff;
  rom[07762] = 16'hffff;
  rom[07763] = 16'hffff;
  rom[07764] = 16'hffff;
  rom[07765] = 16'hffff;
  rom[07766] = 16'hffff;
  rom[07767] = 16'hffff;
  rom[07768] = 16'hffff;
  rom[07769] = 16'hffff;
  rom[07770] = 16'hffff;
  rom[07771] = 16'hffff;
  rom[07772] = 16'hffff;
  rom[07773] = 16'hffff;
  rom[07774] = 16'hffff;
  rom[07775] = 16'hffff;
  rom[07776] = 16'hffff;
  rom[07777] = 16'hffff;
  rom[07778] = 16'hffff;
  rom[07779] = 16'hffff;
  rom[07780] = 16'hffff;
  rom[07781] = 16'hffff;
  rom[07782] = 16'hffff;
  rom[07783] = 16'hffff;
  rom[07784] = 16'hffff;
  rom[07785] = 16'hffff;
  rom[07786] = 16'hffff;
  rom[07787] = 16'hffff;
  rom[07788] = 16'hffff;
  rom[07789] = 16'hffff;
  rom[07790] = 16'hffff;
  rom[07791] = 16'hffff;
  rom[07792] = 16'hffff;
  rom[07793] = 16'hffff;
  rom[07794] = 16'hffff;
  rom[07795] = 16'hffff;
  rom[07796] = 16'hffff;
  rom[07797] = 16'hffff;
  rom[07798] = 16'hffff;
  rom[07799] = 16'hffff;
  rom[07800] = 16'hffff;
  rom[07801] = 16'hffff;
  rom[07802] = 16'hffff;
  rom[07803] = 16'hffff;
  rom[07804] = 16'hffff;
  rom[07805] = 16'hffff;
  rom[07806] = 16'hffff;
  rom[07807] = 16'hffff;
  rom[07808] = 16'hffff;
  rom[07809] = 16'hffff;
  rom[07810] = 16'hffff;
  rom[07811] = 16'hffff;
  rom[07812] = 16'hffff;
  rom[07813] = 16'hffff;
  rom[07814] = 16'hffff;
  rom[07815] = 16'hffff;
  rom[07816] = 16'hffff;
  rom[07817] = 16'hffff;
  rom[07818] = 16'hffff;
  rom[07819] = 16'hffff;
  rom[07820] = 16'hffff;
  rom[07821] = 16'hffff;
  rom[07822] = 16'hffff;
  rom[07823] = 16'hffff;
  rom[07824] = 16'hffff;
  rom[07825] = 16'hffff;
  rom[07826] = 16'hffff;
  rom[07827] = 16'hffff;
  rom[07828] = 16'hffff;
  rom[07829] = 16'hffff;
  rom[07830] = 16'hffff;
  rom[07831] = 16'hffff;
  rom[07832] = 16'hffff;
  rom[07833] = 16'hffff;
  rom[07834] = 16'hffff;
  rom[07835] = 16'hffff;
  rom[07836] = 16'hffff;
  rom[07837] = 16'hffff;
  rom[07838] = 16'hffff;
  rom[07839] = 16'hffff;
  rom[07840] = 16'hffff;
  rom[07841] = 16'hffff;
  rom[07842] = 16'hffff;
  rom[07843] = 16'hffff;
  rom[07844] = 16'hffff;
  rom[07845] = 16'hffff;
  rom[07846] = 16'hffff;
  rom[07847] = 16'hffff;
  rom[07848] = 16'hffff;
  rom[07849] = 16'hffff;
  rom[07850] = 16'hffff;
  rom[07851] = 16'hffff;
  rom[07852] = 16'hffff;
  rom[07853] = 16'hd5f5;
  rom[07854] = 16'h7ae7;
  rom[07855] = 16'hb4cc;
  rom[07856] = 16'hd58f;
  rom[07857] = 16'hc4ed;
  rom[07858] = 16'h4982;
  rom[07859] = 16'h1840;
  rom[07860] = 16'h20c3;
  rom[07861] = 16'h18a3;
  rom[07862] = 16'h18c3;
  rom[07863] = 16'h10a2;
  rom[07864] = 16'h18c2;
  rom[07865] = 16'h18a2;
  rom[07866] = 16'h18a3;
  rom[07867] = 16'h10a3;
  rom[07868] = 16'h18c3;
  rom[07869] = 16'h20e3;
  rom[07870] = 16'h30e1;
  rom[07871] = 16'h93a7;
  rom[07872] = 16'he5cd;
  rom[07873] = 16'hf5c9;
  rom[07874] = 16'hfda8;
  rom[07875] = 16'hfdc8;
  rom[07876] = 16'hfda9;
  rom[07877] = 16'hfdc9;
  rom[07878] = 16'hfde9;
  rom[07879] = 16'hfdc8;
  rom[07880] = 16'hfde9;
  rom[07881] = 16'hf5c8;
  rom[07882] = 16'hfde9;
  rom[07883] = 16'hf5e9;
  rom[07884] = 16'hfe0a;
  rom[07885] = 16'hfde9;
  rom[07886] = 16'hfe0a;
  rom[07887] = 16'hfde9;
  rom[07888] = 16'hfe09;
  rom[07889] = 16'hfde9;
  rom[07890] = 16'hfe0a;
  rom[07891] = 16'hfde9;
  rom[07892] = 16'hfe0a;
  rom[07893] = 16'hfde9;
  rom[07894] = 16'hfe0a;
  rom[07895] = 16'hfde9;
  rom[07896] = 16'hfe0a;
  rom[07897] = 16'hfde9;
  rom[07898] = 16'hfe0a;
  rom[07899] = 16'hfde9;
  rom[07900] = 16'hfe0a;
  rom[07901] = 16'hfde9;
  rom[07902] = 16'hfe0a;
  rom[07903] = 16'hfde9;
  rom[07904] = 16'hfe0a;
  rom[07905] = 16'hfde9;
  rom[07906] = 16'hfdea;
  rom[07907] = 16'hfde9;
  rom[07908] = 16'hfdea;
  rom[07909] = 16'hfde9;
  rom[07910] = 16'hfde9;
  rom[07911] = 16'hfdc8;
  rom[07912] = 16'hfdea;
  rom[07913] = 16'hfdc9;
  rom[07914] = 16'hfdca;
  rom[07915] = 16'hfdc9;
  rom[07916] = 16'hfde9;
  rom[07917] = 16'hf5c8;
  rom[07918] = 16'hfdc8;
  rom[07919] = 16'hfdc8;
  rom[07920] = 16'hfdaa;
  rom[07921] = 16'he54d;
  rom[07922] = 16'h6244;
  rom[07923] = 16'h18a0;
  rom[07924] = 16'h18e3;
  rom[07925] = 16'h08a3;
  rom[07926] = 16'h10e4;
  rom[07927] = 16'h10a2;
  rom[07928] = 16'h20c3;
  rom[07929] = 16'h18a2;
  rom[07930] = 16'h18a3;
  rom[07931] = 16'h1083;
  rom[07932] = 16'h10a4;
  rom[07933] = 16'h18c3;
  rom[07934] = 16'h20c3;
  rom[07935] = 16'h28e0;
  rom[07936] = 16'h9bc8;
  rom[07937] = 16'he56a;
  rom[07938] = 16'hf569;
  rom[07939] = 16'hf54a;
  rom[07940] = 16'hf58d;
  rom[07941] = 16'hcceb;
  rom[07942] = 16'h7b26;
  rom[07943] = 16'he656;
  rom[07944] = 16'hffdf;
  rom[07945] = 16'hffff;
  rom[07946] = 16'hffff;
  rom[07947] = 16'hffff;
  rom[07948] = 16'hffff;
  rom[07949] = 16'hffff;
  rom[07950] = 16'hffff;
  rom[07951] = 16'hffff;
  rom[07952] = 16'hffff;
  rom[07953] = 16'hffff;
  rom[07954] = 16'hffff;
  rom[07955] = 16'hffff;
  rom[07956] = 16'hffff;
  rom[07957] = 16'hffff;
  rom[07958] = 16'hffff;
  rom[07959] = 16'hffff;
  rom[07960] = 16'hffff;
  rom[07961] = 16'hffff;
  rom[07962] = 16'hffff;
  rom[07963] = 16'hffff;
  rom[07964] = 16'hffff;
  rom[07965] = 16'hffff;
  rom[07966] = 16'hffff;
  rom[07967] = 16'hffff;
  rom[07968] = 16'hffff;
  rom[07969] = 16'hffff;
  rom[07970] = 16'hffff;
  rom[07971] = 16'hffff;
  rom[07972] = 16'hffff;
  rom[07973] = 16'hffff;
  rom[07974] = 16'hffff;
  rom[07975] = 16'hffff;
  rom[07976] = 16'hffff;
  rom[07977] = 16'hffff;
  rom[07978] = 16'hffff;
  rom[07979] = 16'hffff;
  rom[07980] = 16'hffff;
  rom[07981] = 16'hffff;
  rom[07982] = 16'hffff;
  rom[07983] = 16'hffff;
  rom[07984] = 16'hffff;
  rom[07985] = 16'hffff;
  rom[07986] = 16'hffff;
  rom[07987] = 16'hffff;
  rom[07988] = 16'hffff;
  rom[07989] = 16'hffff;
  rom[07990] = 16'hffff;
  rom[07991] = 16'hffff;
  rom[07992] = 16'hffff;
  rom[07993] = 16'hffff;
  rom[07994] = 16'hffff;
  rom[07995] = 16'hffff;
  rom[07996] = 16'hffff;
  rom[07997] = 16'hffff;
  rom[07998] = 16'hffff;
  rom[07999] = 16'hffff;
  rom[08000] = 16'hffff;
  rom[08001] = 16'hffff;
  rom[08002] = 16'hffff;
  rom[08003] = 16'hffff;
  rom[08004] = 16'hffff;
  rom[08005] = 16'hffff;
  rom[08006] = 16'hffff;
  rom[08007] = 16'hffff;
  rom[08008] = 16'hffff;
  rom[08009] = 16'hffff;
  rom[08010] = 16'hffff;
  rom[08011] = 16'hffff;
  rom[08012] = 16'hffff;
  rom[08013] = 16'hffff;
  rom[08014] = 16'hffff;
  rom[08015] = 16'hffff;
  rom[08016] = 16'hffff;
  rom[08017] = 16'hffff;
  rom[08018] = 16'hffff;
  rom[08019] = 16'hffff;
  rom[08020] = 16'hffff;
  rom[08021] = 16'hffff;
  rom[08022] = 16'hffff;
  rom[08023] = 16'hffff;
  rom[08024] = 16'hffff;
  rom[08025] = 16'hffff;
  rom[08026] = 16'hffff;
  rom[08027] = 16'hffff;
  rom[08028] = 16'hffff;
  rom[08029] = 16'hffff;
  rom[08030] = 16'hffff;
  rom[08031] = 16'hffff;
  rom[08032] = 16'hffff;
  rom[08033] = 16'hffff;
  rom[08034] = 16'hffff;
  rom[08035] = 16'hffff;
  rom[08036] = 16'hffff;
  rom[08037] = 16'hffff;
  rom[08038] = 16'hffff;
  rom[08039] = 16'hffff;
  rom[08040] = 16'hffff;
  rom[08041] = 16'hffff;
  rom[08042] = 16'hffff;
  rom[08043] = 16'hffff;
  rom[08044] = 16'hffff;
  rom[08045] = 16'hffff;
  rom[08046] = 16'hffff;
  rom[08047] = 16'hffff;
  rom[08048] = 16'hffff;
  rom[08049] = 16'hffff;
  rom[08050] = 16'hffff;
  rom[08051] = 16'hffff;
  rom[08052] = 16'hd636;
  rom[08053] = 16'h7b27;
  rom[08054] = 16'hac49;
  rom[08055] = 16'he5ac;
  rom[08056] = 16'hdd6c;
  rom[08057] = 16'hdd8e;
  rom[08058] = 16'h8307;
  rom[08059] = 16'h30c1;
  rom[08060] = 16'h1881;
  rom[08061] = 16'h10a3;
  rom[08062] = 16'h18c3;
  rom[08063] = 16'h10c3;
  rom[08064] = 16'h10a2;
  rom[08065] = 16'h18a3;
  rom[08066] = 16'h1083;
  rom[08067] = 16'h10a3;
  rom[08068] = 16'h10a2;
  rom[08069] = 16'h1081;
  rom[08070] = 16'h2080;
  rom[08071] = 16'h5a43;
  rom[08072] = 16'hcd0b;
  rom[08073] = 16'hf5cb;
  rom[08074] = 16'hf5a8;
  rom[08075] = 16'hfda9;
  rom[08076] = 16'hfda8;
  rom[08077] = 16'hfdc8;
  rom[08078] = 16'hfde8;
  rom[08079] = 16'hfde9;
  rom[08080] = 16'hf5e9;
  rom[08081] = 16'hf5e9;
  rom[08082] = 16'hfde9;
  rom[08083] = 16'hfde9;
  rom[08084] = 16'hf5e9;
  rom[08085] = 16'hfe09;
  rom[08086] = 16'hfde9;
  rom[08087] = 16'hfe09;
  rom[08088] = 16'hf5e9;
  rom[08089] = 16'hfe09;
  rom[08090] = 16'hfde9;
  rom[08091] = 16'hfe09;
  rom[08092] = 16'hf5e9;
  rom[08093] = 16'hfe09;
  rom[08094] = 16'hfde9;
  rom[08095] = 16'hfe09;
  rom[08096] = 16'hf5e9;
  rom[08097] = 16'hfe09;
  rom[08098] = 16'hfde9;
  rom[08099] = 16'hfe09;
  rom[08100] = 16'hf5e9;
  rom[08101] = 16'hfe09;
  rom[08102] = 16'hfde9;
  rom[08103] = 16'hfe09;
  rom[08104] = 16'hf5e9;
  rom[08105] = 16'hfe09;
  rom[08106] = 16'hfde9;
  rom[08107] = 16'hfe09;
  rom[08108] = 16'hf5e9;
  rom[08109] = 16'hfe09;
  rom[08110] = 16'hfde9;
  rom[08111] = 16'hfde9;
  rom[08112] = 16'hf5c8;
  rom[08113] = 16'hfde8;
  rom[08114] = 16'hfdc9;
  rom[08115] = 16'hfdc9;
  rom[08116] = 16'hf5c9;
  rom[08117] = 16'hfdc8;
  rom[08118] = 16'hfdc8;
  rom[08119] = 16'hf5a8;
  rom[08120] = 16'hedab;
  rom[08121] = 16'habe8;
  rom[08122] = 16'h3100;
  rom[08123] = 16'h18a2;
  rom[08124] = 16'h08c2;
  rom[08125] = 16'h08c3;
  rom[08126] = 16'h10e3;
  rom[08127] = 16'h10c3;
  rom[08128] = 16'h10a2;
  rom[08129] = 16'h18a2;
  rom[08130] = 16'h18a3;
  rom[08131] = 16'h0863;
  rom[08132] = 16'h1084;
  rom[08133] = 16'h18a3;
  rom[08134] = 16'h1860;
  rom[08135] = 16'h6223;
  rom[08136] = 16'hcd29;
  rom[08137] = 16'hf5aa;
  rom[08138] = 16'hf548;
  rom[08139] = 16'hfd6a;
  rom[08140] = 16'hed4a;
  rom[08141] = 16'he56a;
  rom[08142] = 16'ha407;
  rom[08143] = 16'h7b08;
  rom[08144] = 16'heefb;
  rom[08145] = 16'hffff;
  rom[08146] = 16'hffff;
  rom[08147] = 16'hffff;
  rom[08148] = 16'hffff;
  rom[08149] = 16'hffff;
  rom[08150] = 16'hffff;
  rom[08151] = 16'hffff;
  rom[08152] = 16'hffff;
  rom[08153] = 16'hffff;
  rom[08154] = 16'hffff;
  rom[08155] = 16'hffff;
  rom[08156] = 16'hffff;
  rom[08157] = 16'hffff;
  rom[08158] = 16'hffff;
  rom[08159] = 16'hffff;
  rom[08160] = 16'hffff;
  rom[08161] = 16'hffff;
  rom[08162] = 16'hffff;
  rom[08163] = 16'hffff;
  rom[08164] = 16'hffff;
  rom[08165] = 16'hffff;
  rom[08166] = 16'hffff;
  rom[08167] = 16'hffff;
  rom[08168] = 16'hffff;
  rom[08169] = 16'hffff;
  rom[08170] = 16'hffff;
  rom[08171] = 16'hffff;
  rom[08172] = 16'hffff;
  rom[08173] = 16'hffff;
  rom[08174] = 16'hffff;
  rom[08175] = 16'hffff;
  rom[08176] = 16'hffff;
  rom[08177] = 16'hffff;
  rom[08178] = 16'hffff;
  rom[08179] = 16'hffff;
  rom[08180] = 16'hffff;
  rom[08181] = 16'hffff;
  rom[08182] = 16'hffff;
  rom[08183] = 16'hffff;
  rom[08184] = 16'hffff;
  rom[08185] = 16'hffff;
  rom[08186] = 16'hffff;
  rom[08187] = 16'hffff;
  rom[08188] = 16'hffff;
  rom[08189] = 16'hffff;
  rom[08190] = 16'hffff;
  rom[08191] = 16'hffff;
  rom[08192] = 16'hffff;
  rom[08193] = 16'hffff;
  rom[08194] = 16'hffff;
  rom[08195] = 16'hffff;
  rom[08196] = 16'hffff;
  rom[08197] = 16'hffff;
  rom[08198] = 16'hffff;
  rom[08199] = 16'hffff;
  rom[08200] = 16'hffff;
  rom[08201] = 16'hffff;
  rom[08202] = 16'hffff;
  rom[08203] = 16'hffff;
  rom[08204] = 16'hffff;
  rom[08205] = 16'hffff;
  rom[08206] = 16'hffff;
  rom[08207] = 16'hffff;
  rom[08208] = 16'hffff;
  rom[08209] = 16'hffff;
  rom[08210] = 16'hffff;
  rom[08211] = 16'hffff;
  rom[08212] = 16'hffff;
  rom[08213] = 16'hffff;
  rom[08214] = 16'hffff;
  rom[08215] = 16'hffff;
  rom[08216] = 16'hffff;
  rom[08217] = 16'hffff;
  rom[08218] = 16'hffff;
  rom[08219] = 16'hffff;
  rom[08220] = 16'hffff;
  rom[08221] = 16'hffff;
  rom[08222] = 16'hffff;
  rom[08223] = 16'hffff;
  rom[08224] = 16'hffff;
  rom[08225] = 16'hffff;
  rom[08226] = 16'hffff;
  rom[08227] = 16'hffff;
  rom[08228] = 16'hffff;
  rom[08229] = 16'hffff;
  rom[08230] = 16'hffff;
  rom[08231] = 16'hffff;
  rom[08232] = 16'hffff;
  rom[08233] = 16'hffff;
  rom[08234] = 16'hffff;
  rom[08235] = 16'hffff;
  rom[08236] = 16'hffff;
  rom[08237] = 16'hffff;
  rom[08238] = 16'hffff;
  rom[08239] = 16'hffff;
  rom[08240] = 16'hffff;
  rom[08241] = 16'hffff;
  rom[08242] = 16'hffff;
  rom[08243] = 16'hffff;
  rom[08244] = 16'hffff;
  rom[08245] = 16'hffff;
  rom[08246] = 16'hffff;
  rom[08247] = 16'hffff;
  rom[08248] = 16'hffff;
  rom[08249] = 16'hffff;
  rom[08250] = 16'hffff;
  rom[08251] = 16'he6d9;
  rom[08252] = 16'h6285;
  rom[08253] = 16'h9c08;
  rom[08254] = 16'he58c;
  rom[08255] = 16'hf5aa;
  rom[08256] = 16'hf5ab;
  rom[08257] = 16'hdd4b;
  rom[08258] = 16'hbc6b;
  rom[08259] = 16'h4121;
  rom[08260] = 16'h28e1;
  rom[08261] = 16'h10a2;
  rom[08262] = 16'h10c3;
  rom[08263] = 16'h10a3;
  rom[08264] = 16'h10a3;
  rom[08265] = 16'h10a3;
  rom[08266] = 16'h10a3;
  rom[08267] = 16'h10a3;
  rom[08268] = 16'h10c3;
  rom[08269] = 16'h1082;
  rom[08270] = 16'h20c2;
  rom[08271] = 16'h28e0;
  rom[08272] = 16'h9ba8;
  rom[08273] = 16'he56b;
  rom[08274] = 16'hfdeb;
  rom[08275] = 16'hfda9;
  rom[08276] = 16'hfde9;
  rom[08277] = 16'hfda7;
  rom[08278] = 16'hfde9;
  rom[08279] = 16'hfdc9;
  rom[08280] = 16'hfdea;
  rom[08281] = 16'hf5c9;
  rom[08282] = 16'hfe0a;
  rom[08283] = 16'hfde9;
  rom[08284] = 16'hfe0a;
  rom[08285] = 16'hfde9;
  rom[08286] = 16'hfe0a;
  rom[08287] = 16'hfde9;
  rom[08288] = 16'hfe0a;
  rom[08289] = 16'hfde9;
  rom[08290] = 16'hfe0a;
  rom[08291] = 16'hfde9;
  rom[08292] = 16'hfe0a;
  rom[08293] = 16'hfde9;
  rom[08294] = 16'hfe0a;
  rom[08295] = 16'hfde9;
  rom[08296] = 16'hfe0a;
  rom[08297] = 16'hfde9;
  rom[08298] = 16'hfe0a;
  rom[08299] = 16'hfde9;
  rom[08300] = 16'hfe0a;
  rom[08301] = 16'hfde9;
  rom[08302] = 16'hfe0a;
  rom[08303] = 16'hfde9;
  rom[08304] = 16'hfe0a;
  rom[08305] = 16'hfde9;
  rom[08306] = 16'hfe0a;
  rom[08307] = 16'hfde9;
  rom[08308] = 16'hfe0a;
  rom[08309] = 16'hfde9;
  rom[08310] = 16'hfe0a;
  rom[08311] = 16'hfde9;
  rom[08312] = 16'hfe09;
  rom[08313] = 16'hfdc7;
  rom[08314] = 16'hfde9;
  rom[08315] = 16'hfdc9;
  rom[08316] = 16'hfdea;
  rom[08317] = 16'hfde9;
  rom[08318] = 16'hfde9;
  rom[08319] = 16'hf5e9;
  rom[08320] = 16'he58c;
  rom[08321] = 16'h7ae6;
  rom[08322] = 16'h28a1;
  rom[08323] = 16'h18a2;
  rom[08324] = 16'h08a2;
  rom[08325] = 16'h08c2;
  rom[08326] = 16'h10e3;
  rom[08327] = 16'h08c2;
  rom[08328] = 16'h10c2;
  rom[08329] = 16'h10a2;
  rom[08330] = 16'h18c3;
  rom[08331] = 16'h10a3;
  rom[08332] = 16'h18c5;
  rom[08333] = 16'h20a3;
  rom[08334] = 16'h38e1;
  rom[08335] = 16'h9365;
  rom[08336] = 16'hf60a;
  rom[08337] = 16'hf5a9;
  rom[08338] = 16'hfd28;
  rom[08339] = 16'hfd69;
  rom[08340] = 16'hf549;
  rom[08341] = 16'hf5c9;
  rom[08342] = 16'hdd6b;
  rom[08343] = 16'h8305;
  rom[08344] = 16'hbcf3;
  rom[08345] = 16'hffff;
  rom[08346] = 16'hffff;
  rom[08347] = 16'hffff;
  rom[08348] = 16'hffff;
  rom[08349] = 16'hffff;
  rom[08350] = 16'hffff;
  rom[08351] = 16'hffff;
  rom[08352] = 16'hffff;
  rom[08353] = 16'hffff;
  rom[08354] = 16'hffff;
  rom[08355] = 16'hffff;
  rom[08356] = 16'hffff;
  rom[08357] = 16'hffff;
  rom[08358] = 16'hffff;
  rom[08359] = 16'hffff;
  rom[08360] = 16'hffff;
  rom[08361] = 16'hffff;
  rom[08362] = 16'hffff;
  rom[08363] = 16'hffff;
  rom[08364] = 16'hffff;
  rom[08365] = 16'hffff;
  rom[08366] = 16'hffff;
  rom[08367] = 16'hffff;
  rom[08368] = 16'hffff;
  rom[08369] = 16'hffff;
  rom[08370] = 16'hffff;
  rom[08371] = 16'hffff;
  rom[08372] = 16'hffff;
  rom[08373] = 16'hffff;
  rom[08374] = 16'hffff;
  rom[08375] = 16'hffff;
  rom[08376] = 16'hffff;
  rom[08377] = 16'hffff;
  rom[08378] = 16'hffff;
  rom[08379] = 16'hffff;
  rom[08380] = 16'hffff;
  rom[08381] = 16'hffff;
  rom[08382] = 16'hffff;
  rom[08383] = 16'hffff;
  rom[08384] = 16'hffff;
  rom[08385] = 16'hffff;
  rom[08386] = 16'hffff;
  rom[08387] = 16'hffff;
  rom[08388] = 16'hffff;
  rom[08389] = 16'hffff;
  rom[08390] = 16'hffff;
  rom[08391] = 16'hffff;
  rom[08392] = 16'hffff;
  rom[08393] = 16'hffff;
  rom[08394] = 16'hffff;
  rom[08395] = 16'hffff;
  rom[08396] = 16'hffff;
  rom[08397] = 16'hffff;
  rom[08398] = 16'hffff;
  rom[08399] = 16'hffff;
  rom[08400] = 16'hffff;
  rom[08401] = 16'hffff;
  rom[08402] = 16'hffff;
  rom[08403] = 16'hffff;
  rom[08404] = 16'hffff;
  rom[08405] = 16'hffff;
  rom[08406] = 16'hffff;
  rom[08407] = 16'hffff;
  rom[08408] = 16'hffff;
  rom[08409] = 16'hffff;
  rom[08410] = 16'hffff;
  rom[08411] = 16'hffff;
  rom[08412] = 16'hffff;
  rom[08413] = 16'hffff;
  rom[08414] = 16'hffff;
  rom[08415] = 16'hffff;
  rom[08416] = 16'hffff;
  rom[08417] = 16'hffff;
  rom[08418] = 16'hffff;
  rom[08419] = 16'hffff;
  rom[08420] = 16'hffff;
  rom[08421] = 16'hffff;
  rom[08422] = 16'hffff;
  rom[08423] = 16'hffff;
  rom[08424] = 16'hffff;
  rom[08425] = 16'hffff;
  rom[08426] = 16'hffff;
  rom[08427] = 16'hffff;
  rom[08428] = 16'hffff;
  rom[08429] = 16'hffff;
  rom[08430] = 16'hffff;
  rom[08431] = 16'hffff;
  rom[08432] = 16'hffff;
  rom[08433] = 16'hffff;
  rom[08434] = 16'hffff;
  rom[08435] = 16'hffff;
  rom[08436] = 16'hffff;
  rom[08437] = 16'hffff;
  rom[08438] = 16'hffff;
  rom[08439] = 16'hffff;
  rom[08440] = 16'hffff;
  rom[08441] = 16'hffff;
  rom[08442] = 16'hffff;
  rom[08443] = 16'hffff;
  rom[08444] = 16'hffff;
  rom[08445] = 16'hffff;
  rom[08446] = 16'hffdf;
  rom[08447] = 16'hffdf;
  rom[08448] = 16'hffff;
  rom[08449] = 16'hffff;
  rom[08450] = 16'hffbc;
  rom[08451] = 16'h7b69;
  rom[08452] = 16'ha428;
  rom[08453] = 16'hdd8b;
  rom[08454] = 16'hedaa;
  rom[08455] = 16'hfd88;
  rom[08456] = 16'hf568;
  rom[08457] = 16'hf56b;
  rom[08458] = 16'he54c;
  rom[08459] = 16'h7ac5;
  rom[08460] = 16'h28c0;
  rom[08461] = 16'h20c1;
  rom[08462] = 16'h10a2;
  rom[08463] = 16'h10a3;
  rom[08464] = 16'h10a3;
  rom[08465] = 16'h10a3;
  rom[08466] = 16'h10a3;
  rom[08467] = 16'h10c3;
  rom[08468] = 16'h10a3;
  rom[08469] = 16'h10a3;
  rom[08470] = 16'h10c2;
  rom[08471] = 16'h18a0;
  rom[08472] = 16'h5a24;
  rom[08473] = 16'hcd2d;
  rom[08474] = 16'hedab;
  rom[08475] = 16'hfdea;
  rom[08476] = 16'hfda7;
  rom[08477] = 16'hfdc7;
  rom[08478] = 16'hfde8;
  rom[08479] = 16'hf5c9;
  rom[08480] = 16'hf5e9;
  rom[08481] = 16'hf5e9;
  rom[08482] = 16'hf5c9;
  rom[08483] = 16'hfde9;
  rom[08484] = 16'hf5e9;
  rom[08485] = 16'hfe09;
  rom[08486] = 16'hf5e9;
  rom[08487] = 16'hfe09;
  rom[08488] = 16'hfde9;
  rom[08489] = 16'hfe09;
  rom[08490] = 16'hf5e9;
  rom[08491] = 16'hfe09;
  rom[08492] = 16'hfde9;
  rom[08493] = 16'hfe09;
  rom[08494] = 16'hf5e9;
  rom[08495] = 16'hfe09;
  rom[08496] = 16'hfde9;
  rom[08497] = 16'hfe09;
  rom[08498] = 16'hf5e9;
  rom[08499] = 16'hfe09;
  rom[08500] = 16'hfde9;
  rom[08501] = 16'hfe09;
  rom[08502] = 16'hf5e9;
  rom[08503] = 16'hfe09;
  rom[08504] = 16'hfde9;
  rom[08505] = 16'hfe09;
  rom[08506] = 16'hf5e9;
  rom[08507] = 16'hfe09;
  rom[08508] = 16'hfde9;
  rom[08509] = 16'hfe09;
  rom[08510] = 16'hf5c8;
  rom[08511] = 16'hfde9;
  rom[08512] = 16'hfdc8;
  rom[08513] = 16'hfde8;
  rom[08514] = 16'hf5c8;
  rom[08515] = 16'hfde9;
  rom[08516] = 16'hfdc9;
  rom[08517] = 16'hfde9;
  rom[08518] = 16'hedc9;
  rom[08519] = 16'hf62c;
  rom[08520] = 16'hbceb;
  rom[08521] = 16'h3942;
  rom[08522] = 16'h1881;
  rom[08523] = 16'h18a3;
  rom[08524] = 16'h08a2;
  rom[08525] = 16'h10e2;
  rom[08526] = 16'h10c2;
  rom[08527] = 16'h10a3;
  rom[08528] = 16'h10a2;
  rom[08529] = 16'h10a2;
  rom[08530] = 16'h10a2;
  rom[08531] = 16'h18c3;
  rom[08532] = 16'h1062;
  rom[08533] = 16'h28a1;
  rom[08534] = 16'h59e2;
  rom[08535] = 16'hd50a;
  rom[08536] = 16'hedc8;
  rom[08537] = 16'hfd88;
  rom[08538] = 16'hf528;
  rom[08539] = 16'hfd69;
  rom[08540] = 16'hf569;
  rom[08541] = 16'hf589;
  rom[08542] = 16'he56a;
  rom[08543] = 16'hccec;
  rom[08544] = 16'h7ac7;
  rom[08545] = 16'hf6fb;
  rom[08546] = 16'hffbf;
  rom[08547] = 16'hffff;
  rom[08548] = 16'hffff;
  rom[08549] = 16'hffff;
  rom[08550] = 16'hffff;
  rom[08551] = 16'hffff;
  rom[08552] = 16'hffff;
  rom[08553] = 16'hffff;
  rom[08554] = 16'hffff;
  rom[08555] = 16'hffff;
  rom[08556] = 16'hffff;
  rom[08557] = 16'hffff;
  rom[08558] = 16'hffff;
  rom[08559] = 16'hffff;
  rom[08560] = 16'hffff;
  rom[08561] = 16'hffff;
  rom[08562] = 16'hffff;
  rom[08563] = 16'hffff;
  rom[08564] = 16'hffff;
  rom[08565] = 16'hffff;
  rom[08566] = 16'hffff;
  rom[08567] = 16'hffff;
  rom[08568] = 16'hffff;
  rom[08569] = 16'hffff;
  rom[08570] = 16'hffff;
  rom[08571] = 16'hffff;
  rom[08572] = 16'hffff;
  rom[08573] = 16'hffff;
  rom[08574] = 16'hffff;
  rom[08575] = 16'hffff;
  rom[08576] = 16'hffff;
  rom[08577] = 16'hffff;
  rom[08578] = 16'hffff;
  rom[08579] = 16'hffff;
  rom[08580] = 16'hffff;
  rom[08581] = 16'hffff;
  rom[08582] = 16'hffff;
  rom[08583] = 16'hffff;
  rom[08584] = 16'hffff;
  rom[08585] = 16'hffff;
  rom[08586] = 16'hffff;
  rom[08587] = 16'hffff;
  rom[08588] = 16'hffff;
  rom[08589] = 16'hffff;
  rom[08590] = 16'hffff;
  rom[08591] = 16'hffff;
  rom[08592] = 16'hffff;
  rom[08593] = 16'hffff;
  rom[08594] = 16'hffff;
  rom[08595] = 16'hffff;
  rom[08596] = 16'hffff;
  rom[08597] = 16'hffff;
  rom[08598] = 16'hffff;
  rom[08599] = 16'hffff;
  rom[08600] = 16'hffff;
  rom[08601] = 16'hffff;
  rom[08602] = 16'hffff;
  rom[08603] = 16'hffff;
  rom[08604] = 16'hffff;
  rom[08605] = 16'hffff;
  rom[08606] = 16'hffff;
  rom[08607] = 16'hffff;
  rom[08608] = 16'hffff;
  rom[08609] = 16'hffff;
  rom[08610] = 16'hffff;
  rom[08611] = 16'hffff;
  rom[08612] = 16'hffff;
  rom[08613] = 16'hffff;
  rom[08614] = 16'hffff;
  rom[08615] = 16'hffff;
  rom[08616] = 16'hffff;
  rom[08617] = 16'hffff;
  rom[08618] = 16'hffff;
  rom[08619] = 16'hffff;
  rom[08620] = 16'hffff;
  rom[08621] = 16'hffff;
  rom[08622] = 16'hffff;
  rom[08623] = 16'hffff;
  rom[08624] = 16'hffff;
  rom[08625] = 16'hffff;
  rom[08626] = 16'hffff;
  rom[08627] = 16'hffff;
  rom[08628] = 16'hffff;
  rom[08629] = 16'hffff;
  rom[08630] = 16'hffff;
  rom[08631] = 16'hffff;
  rom[08632] = 16'hffff;
  rom[08633] = 16'hffff;
  rom[08634] = 16'hffff;
  rom[08635] = 16'hffff;
  rom[08636] = 16'hffff;
  rom[08637] = 16'hffff;
  rom[08638] = 16'hffff;
  rom[08639] = 16'hffff;
  rom[08640] = 16'hffff;
  rom[08641] = 16'hffff;
  rom[08642] = 16'hffff;
  rom[08643] = 16'hffff;
  rom[08644] = 16'hffff;
  rom[08645] = 16'hfffe;
  rom[08646] = 16'hffff;
  rom[08647] = 16'hffff;
  rom[08648] = 16'hff9e;
  rom[08649] = 16'hff9d;
  rom[08650] = 16'h8b8b;
  rom[08651] = 16'h8325;
  rom[08652] = 16'hdd6c;
  rom[08653] = 16'hedaa;
  rom[08654] = 16'hfda8;
  rom[08655] = 16'hf526;
  rom[08656] = 16'hfd69;
  rom[08657] = 16'hfd4a;
  rom[08658] = 16'hf58c;
  rom[08659] = 16'hc4eb;
  rom[08660] = 16'h49a1;
  rom[08661] = 16'h20c1;
  rom[08662] = 16'h18a1;
  rom[08663] = 16'h18a2;
  rom[08664] = 16'h18a3;
  rom[08665] = 16'h10a3;
  rom[08666] = 16'h10c3;
  rom[08667] = 16'h10c3;
  rom[08668] = 16'h10c3;
  rom[08669] = 16'h10a3;
  rom[08670] = 16'h10c3;
  rom[08671] = 16'h10c2;
  rom[08672] = 16'h28c1;
  rom[08673] = 16'ha40a;
  rom[08674] = 16'he58d;
  rom[08675] = 16'hfdea;
  rom[08676] = 16'hfde8;
  rom[08677] = 16'hfe08;
  rom[08678] = 16'hfdc8;
  rom[08679] = 16'hf5c8;
  rom[08680] = 16'hfe0a;
  rom[08681] = 16'hfde9;
  rom[08682] = 16'hfde9;
  rom[08683] = 16'hfde9;
  rom[08684] = 16'hfe09;
  rom[08685] = 16'hfde8;
  rom[08686] = 16'hfe0a;
  rom[08687] = 16'hfde9;
  rom[08688] = 16'hfe0a;
  rom[08689] = 16'hfde9;
  rom[08690] = 16'hfe0a;
  rom[08691] = 16'hfde9;
  rom[08692] = 16'hfe0a;
  rom[08693] = 16'hfde9;
  rom[08694] = 16'hfe0a;
  rom[08695] = 16'hfde9;
  rom[08696] = 16'hfe0a;
  rom[08697] = 16'hfde9;
  rom[08698] = 16'hfe0a;
  rom[08699] = 16'hfde9;
  rom[08700] = 16'hfe0a;
  rom[08701] = 16'hfe09;
  rom[08702] = 16'hfe2a;
  rom[08703] = 16'hfe09;
  rom[08704] = 16'hfe0a;
  rom[08705] = 16'hfde9;
  rom[08706] = 16'hfe0a;
  rom[08707] = 16'hfde9;
  rom[08708] = 16'hfe0a;
  rom[08709] = 16'hfde9;
  rom[08710] = 16'hfe09;
  rom[08711] = 16'hfdc8;
  rom[08712] = 16'hfe09;
  rom[08713] = 16'hf5e9;
  rom[08714] = 16'hfe2a;
  rom[08715] = 16'hf5c8;
  rom[08716] = 16'hfde9;
  rom[08717] = 16'hfde9;
  rom[08718] = 16'hedca;
  rom[08719] = 16'hee0e;
  rom[08720] = 16'h72c6;
  rom[08721] = 16'h20c1;
  rom[08722] = 16'h18c2;
  rom[08723] = 16'h10c3;
  rom[08724] = 16'h10c2;
  rom[08725] = 16'h10a1;
  rom[08726] = 16'h10c2;
  rom[08727] = 16'h10a3;
  rom[08728] = 16'h18a3;
  rom[08729] = 16'h18a2;
  rom[08730] = 16'h10a1;
  rom[08731] = 16'h10a2;
  rom[08732] = 16'h20a2;
  rom[08733] = 16'h28a0;
  rom[08734] = 16'hbc6a;
  rom[08735] = 16'he56a;
  rom[08736] = 16'hf5a9;
  rom[08737] = 16'hfd88;
  rom[08738] = 16'hfd88;
  rom[08739] = 16'hf548;
  rom[08740] = 16'hf569;
  rom[08741] = 16'hf548;
  rom[08742] = 16'hf56a;
  rom[08743] = 16'hed6c;
  rom[08744] = 16'ha389;
  rom[08745] = 16'ha3ee;
  rom[08746] = 16'hffbe;
  rom[08747] = 16'hffff;
  rom[08748] = 16'hffff;
  rom[08749] = 16'hffff;
  rom[08750] = 16'hffff;
  rom[08751] = 16'hffff;
  rom[08752] = 16'hffff;
  rom[08753] = 16'hffff;
  rom[08754] = 16'hffff;
  rom[08755] = 16'hffff;
  rom[08756] = 16'hffff;
  rom[08757] = 16'hffff;
  rom[08758] = 16'hffff;
  rom[08759] = 16'hffff;
  rom[08760] = 16'hffff;
  rom[08761] = 16'hffff;
  rom[08762] = 16'hffff;
  rom[08763] = 16'hffff;
  rom[08764] = 16'hffff;
  rom[08765] = 16'hffff;
  rom[08766] = 16'hffff;
  rom[08767] = 16'hffff;
  rom[08768] = 16'hffff;
  rom[08769] = 16'hffff;
  rom[08770] = 16'hffff;
  rom[08771] = 16'hffff;
  rom[08772] = 16'hffff;
  rom[08773] = 16'hffff;
  rom[08774] = 16'hffff;
  rom[08775] = 16'hffff;
  rom[08776] = 16'hffff;
  rom[08777] = 16'hffff;
  rom[08778] = 16'hffff;
  rom[08779] = 16'hffff;
  rom[08780] = 16'hffff;
  rom[08781] = 16'hffff;
  rom[08782] = 16'hffff;
  rom[08783] = 16'hffff;
  rom[08784] = 16'hffff;
  rom[08785] = 16'hffff;
  rom[08786] = 16'hffff;
  rom[08787] = 16'hffff;
  rom[08788] = 16'hffff;
  rom[08789] = 16'hffff;
  rom[08790] = 16'hffff;
  rom[08791] = 16'hffff;
  rom[08792] = 16'hffff;
  rom[08793] = 16'hffff;
  rom[08794] = 16'hffff;
  rom[08795] = 16'hffff;
  rom[08796] = 16'hffff;
  rom[08797] = 16'hffff;
  rom[08798] = 16'hffff;
  rom[08799] = 16'hffff;
  rom[08800] = 16'hffff;
  rom[08801] = 16'hffff;
  rom[08802] = 16'hffff;
  rom[08803] = 16'hffff;
  rom[08804] = 16'hffff;
  rom[08805] = 16'hffff;
  rom[08806] = 16'hffff;
  rom[08807] = 16'hffff;
  rom[08808] = 16'hffff;
  rom[08809] = 16'hffff;
  rom[08810] = 16'hffff;
  rom[08811] = 16'hffff;
  rom[08812] = 16'hffff;
  rom[08813] = 16'hffff;
  rom[08814] = 16'hffff;
  rom[08815] = 16'hffff;
  rom[08816] = 16'hffff;
  rom[08817] = 16'hffff;
  rom[08818] = 16'hffff;
  rom[08819] = 16'hffff;
  rom[08820] = 16'hffff;
  rom[08821] = 16'hffff;
  rom[08822] = 16'hffff;
  rom[08823] = 16'hffff;
  rom[08824] = 16'hffff;
  rom[08825] = 16'hffff;
  rom[08826] = 16'hffff;
  rom[08827] = 16'hffff;
  rom[08828] = 16'hffff;
  rom[08829] = 16'hffff;
  rom[08830] = 16'hffff;
  rom[08831] = 16'hffff;
  rom[08832] = 16'hffff;
  rom[08833] = 16'hffff;
  rom[08834] = 16'hffff;
  rom[08835] = 16'hffff;
  rom[08836] = 16'hffff;
  rom[08837] = 16'hffff;
  rom[08838] = 16'hffff;
  rom[08839] = 16'hffff;
  rom[08840] = 16'hffff;
  rom[08841] = 16'hffff;
  rom[08842] = 16'hffff;
  rom[08843] = 16'hffff;
  rom[08844] = 16'hffff;
  rom[08845] = 16'hffff;
  rom[08846] = 16'hffff;
  rom[08847] = 16'hffff;
  rom[08848] = 16'hffbe;
  rom[08849] = 16'hbcf1;
  rom[08850] = 16'h6a44;
  rom[08851] = 16'hdd4d;
  rom[08852] = 16'he56a;
  rom[08853] = 16'hf569;
  rom[08854] = 16'hfd68;
  rom[08855] = 16'hfd89;
  rom[08856] = 16'hfd27;
  rom[08857] = 16'hfd69;
  rom[08858] = 16'hf56a;
  rom[08859] = 16'hedad;
  rom[08860] = 16'h8366;
  rom[08861] = 16'h3121;
  rom[08862] = 16'h18a0;
  rom[08863] = 16'h18c2;
  rom[08864] = 16'h18a2;
  rom[08865] = 16'h10a2;
  rom[08866] = 16'h10a2;
  rom[08867] = 16'h10c2;
  rom[08868] = 16'h10a3;
  rom[08869] = 16'h10c3;
  rom[08870] = 16'h10a3;
  rom[08871] = 16'h18e3;
  rom[08872] = 16'h1860;
  rom[08873] = 16'h6244;
  rom[08874] = 16'hd56d;
  rom[08875] = 16'hf5eb;
  rom[08876] = 16'hf5a7;
  rom[08877] = 16'hfe08;
  rom[08878] = 16'hfdc8;
  rom[08879] = 16'hf5c9;
  rom[08880] = 16'hf5e9;
  rom[08881] = 16'hfe09;
  rom[08882] = 16'hf5e9;
  rom[08883] = 16'hfe29;
  rom[08884] = 16'hf5e8;
  rom[08885] = 16'hfe08;
  rom[08886] = 16'hfde8;
  rom[08887] = 16'hfe09;
  rom[08888] = 16'hf608;
  rom[08889] = 16'hfe29;
  rom[08890] = 16'hfe09;
  rom[08891] = 16'hfe29;
  rom[08892] = 16'hf609;
  rom[08893] = 16'hfe29;
  rom[08894] = 16'hfe09;
  rom[08895] = 16'hfe29;
  rom[08896] = 16'hf609;
  rom[08897] = 16'hfe29;
  rom[08898] = 16'hfe09;
  rom[08899] = 16'hfe29;
  rom[08900] = 16'hf609;
  rom[08901] = 16'hfe29;
  rom[08902] = 16'hfe09;
  rom[08903] = 16'hfe29;
  rom[08904] = 16'hf609;
  rom[08905] = 16'hfe29;
  rom[08906] = 16'hfe09;
  rom[08907] = 16'hfe09;
  rom[08908] = 16'hf5e9;
  rom[08909] = 16'hfe09;
  rom[08910] = 16'hfde9;
  rom[08911] = 16'hfe09;
  rom[08912] = 16'hf5e9;
  rom[08913] = 16'hf609;
  rom[08914] = 16'hf5c8;
  rom[08915] = 16'hfde8;
  rom[08916] = 16'hf5e8;
  rom[08917] = 16'hf5e9;
  rom[08918] = 16'he60c;
  rom[08919] = 16'hc52d;
  rom[08920] = 16'h3982;
  rom[08921] = 16'h18c2;
  rom[08922] = 16'h0882;
  rom[08923] = 16'h10a3;
  rom[08924] = 16'h18c2;
  rom[08925] = 16'h10a2;
  rom[08926] = 16'h18c2;
  rom[08927] = 16'h10c3;
  rom[08928] = 16'h10a2;
  rom[08929] = 16'h18c2;
  rom[08930] = 16'h18c1;
  rom[08931] = 16'h18a2;
  rom[08932] = 16'h28c1;
  rom[08933] = 16'h7ac7;
  rom[08934] = 16'hdd6c;
  rom[08935] = 16'hf5ab;
  rom[08936] = 16'hf548;
  rom[08937] = 16'hfd68;
  rom[08938] = 16'hfd47;
  rom[08939] = 16'hfd68;
  rom[08940] = 16'hf568;
  rom[08941] = 16'hfd49;
  rom[08942] = 16'hf569;
  rom[08943] = 16'hed2a;
  rom[08944] = 16'hd50c;
  rom[08945] = 16'h5982;
  rom[08946] = 16'hde78;
  rom[08947] = 16'hffff;
  rom[08948] = 16'hffff;
  rom[08949] = 16'hffff;
  rom[08950] = 16'hffff;
  rom[08951] = 16'hffdf;
  rom[08952] = 16'hffff;
  rom[08953] = 16'hffff;
  rom[08954] = 16'hffff;
  rom[08955] = 16'hffff;
  rom[08956] = 16'hffff;
  rom[08957] = 16'hffff;
  rom[08958] = 16'hffff;
  rom[08959] = 16'hffff;
  rom[08960] = 16'hffff;
  rom[08961] = 16'hffff;
  rom[08962] = 16'hffff;
  rom[08963] = 16'hffff;
  rom[08964] = 16'hffff;
  rom[08965] = 16'hffff;
  rom[08966] = 16'hffff;
  rom[08967] = 16'hffff;
  rom[08968] = 16'hffff;
  rom[08969] = 16'hffff;
  rom[08970] = 16'hffff;
  rom[08971] = 16'hffff;
  rom[08972] = 16'hffff;
  rom[08973] = 16'hffff;
  rom[08974] = 16'hffff;
  rom[08975] = 16'hffff;
  rom[08976] = 16'hffff;
  rom[08977] = 16'hffff;
  rom[08978] = 16'hffff;
  rom[08979] = 16'hffff;
  rom[08980] = 16'hffff;
  rom[08981] = 16'hffff;
  rom[08982] = 16'hffff;
  rom[08983] = 16'hffff;
  rom[08984] = 16'hffff;
  rom[08985] = 16'hffff;
  rom[08986] = 16'hffff;
  rom[08987] = 16'hffff;
  rom[08988] = 16'hffff;
  rom[08989] = 16'hffff;
  rom[08990] = 16'hffff;
  rom[08991] = 16'hffff;
  rom[08992] = 16'hffff;
  rom[08993] = 16'hffff;
  rom[08994] = 16'hffff;
  rom[08995] = 16'hffff;
  rom[08996] = 16'hffff;
  rom[08997] = 16'hffff;
  rom[08998] = 16'hffff;
  rom[08999] = 16'hffff;
  rom[09000] = 16'hffff;
  rom[09001] = 16'hffff;
  rom[09002] = 16'hffff;
  rom[09003] = 16'hffff;
  rom[09004] = 16'hffff;
  rom[09005] = 16'hffff;
  rom[09006] = 16'hffff;
  rom[09007] = 16'hffff;
  rom[09008] = 16'hffff;
  rom[09009] = 16'hffff;
  rom[09010] = 16'hffff;
  rom[09011] = 16'hffff;
  rom[09012] = 16'hffff;
  rom[09013] = 16'hffff;
  rom[09014] = 16'hffff;
  rom[09015] = 16'hffff;
  rom[09016] = 16'hffff;
  rom[09017] = 16'hffff;
  rom[09018] = 16'hffff;
  rom[09019] = 16'hffff;
  rom[09020] = 16'hffff;
  rom[09021] = 16'hffff;
  rom[09022] = 16'hffff;
  rom[09023] = 16'hffff;
  rom[09024] = 16'hffff;
  rom[09025] = 16'hffff;
  rom[09026] = 16'hffff;
  rom[09027] = 16'hffff;
  rom[09028] = 16'hffff;
  rom[09029] = 16'hffff;
  rom[09030] = 16'hffff;
  rom[09031] = 16'hffff;
  rom[09032] = 16'hffff;
  rom[09033] = 16'hffff;
  rom[09034] = 16'hffff;
  rom[09035] = 16'hffff;
  rom[09036] = 16'hffff;
  rom[09037] = 16'hffff;
  rom[09038] = 16'hffff;
  rom[09039] = 16'hffff;
  rom[09040] = 16'hffff;
  rom[09041] = 16'hffff;
  rom[09042] = 16'hffff;
  rom[09043] = 16'hffff;
  rom[09044] = 16'hffff;
  rom[09045] = 16'hffff;
  rom[09046] = 16'hffff;
  rom[09047] = 16'hffdf;
  rom[09048] = 16'hf6b9;
  rom[09049] = 16'h7ae6;
  rom[09050] = 16'hdd8d;
  rom[09051] = 16'he549;
  rom[09052] = 16'hfdaa;
  rom[09053] = 16'hfd49;
  rom[09054] = 16'hfd6a;
  rom[09055] = 16'hfd49;
  rom[09056] = 16'hfd47;
  rom[09057] = 16'hfd88;
  rom[09058] = 16'hfdca;
  rom[09059] = 16'he58b;
  rom[09060] = 16'hd56e;
  rom[09061] = 16'h5a23;
  rom[09062] = 16'h18a1;
  rom[09063] = 16'h18e2;
  rom[09064] = 16'h18a2;
  rom[09065] = 16'h1082;
  rom[09066] = 16'h18c3;
  rom[09067] = 16'h18a2;
  rom[09068] = 16'h18c2;
  rom[09069] = 16'h10a3;
  rom[09070] = 16'h1083;
  rom[09071] = 16'h1083;
  rom[09072] = 16'h20c3;
  rom[09073] = 16'h20a0;
  rom[09074] = 16'hac6a;
  rom[09075] = 16'he5cc;
  rom[09076] = 16'hfe0a;
  rom[09077] = 16'hfde8;
  rom[09078] = 16'hfe09;
  rom[09079] = 16'hfdc8;
  rom[09080] = 16'hfde9;
  rom[09081] = 16'hfde9;
  rom[09082] = 16'hfdc9;
  rom[09083] = 16'hfe2a;
  rom[09084] = 16'hfde9;
  rom[09085] = 16'hfe08;
  rom[09086] = 16'hfe29;
  rom[09087] = 16'hf628;
  rom[09088] = 16'hf629;
  rom[09089] = 16'hf629;
  rom[09090] = 16'hfe2a;
  rom[09091] = 16'hfe29;
  rom[09092] = 16'hfe2a;
  rom[09093] = 16'hfe09;
  rom[09094] = 16'hfe2b;
  rom[09095] = 16'hfe09;
  rom[09096] = 16'hfe2a;
  rom[09097] = 16'hfe29;
  rom[09098] = 16'hfe2a;
  rom[09099] = 16'hfe2a;
  rom[09100] = 16'hfe2a;
  rom[09101] = 16'hfe2a;
  rom[09102] = 16'hfe2a;
  rom[09103] = 16'hfe09;
  rom[09104] = 16'hfe2a;
  rom[09105] = 16'hfe2a;
  rom[09106] = 16'hfdea;
  rom[09107] = 16'hfde9;
  rom[09108] = 16'hfe09;
  rom[09109] = 16'hfe09;
  rom[09110] = 16'hfe29;
  rom[09111] = 16'hf609;
  rom[09112] = 16'hfe29;
  rom[09113] = 16'hf609;
  rom[09114] = 16'hf5c7;
  rom[09115] = 16'hf607;
  rom[09116] = 16'hf627;
  rom[09117] = 16'hede9;
  rom[09118] = 16'heded;
  rom[09119] = 16'h7ae6;
  rom[09120] = 16'h20a1;
  rom[09121] = 16'h10a2;
  rom[09122] = 16'h18c3;
  rom[09123] = 16'h10a2;
  rom[09124] = 16'h18c3;
  rom[09125] = 16'h18c3;
  rom[09126] = 16'h18a2;
  rom[09127] = 16'h18c2;
  rom[09128] = 16'h1883;
  rom[09129] = 16'h18a3;
  rom[09130] = 16'h18a2;
  rom[09131] = 16'h20c1;
  rom[09132] = 16'h4983;
  rom[09133] = 16'hcd4d;
  rom[09134] = 16'hf5ec;
  rom[09135] = 16'hed28;
  rom[09136] = 16'hfdaa;
  rom[09137] = 16'hfd69;
  rom[09138] = 16'hfd89;
  rom[09139] = 16'hfd68;
  rom[09140] = 16'hfd69;
  rom[09141] = 16'hfd49;
  rom[09142] = 16'hfd68;
  rom[09143] = 16'hf568;
  rom[09144] = 16'hed8b;
  rom[09145] = 16'ha3c8;
  rom[09146] = 16'h8b8b;
  rom[09147] = 16'hffbe;
  rom[09148] = 16'hffff;
  rom[09149] = 16'hffff;
  rom[09150] = 16'hf75e;
  rom[09151] = 16'hbdb6;
  rom[09152] = 16'hffbf;
  rom[09153] = 16'hffff;
  rom[09154] = 16'hffff;
  rom[09155] = 16'hffff;
  rom[09156] = 16'hffff;
  rom[09157] = 16'hffff;
  rom[09158] = 16'hffff;
  rom[09159] = 16'hffff;
  rom[09160] = 16'hffff;
  rom[09161] = 16'hffff;
  rom[09162] = 16'hffff;
  rom[09163] = 16'hffff;
  rom[09164] = 16'hffff;
  rom[09165] = 16'hffff;
  rom[09166] = 16'hffff;
  rom[09167] = 16'hffff;
  rom[09168] = 16'hffff;
  rom[09169] = 16'hffff;
  rom[09170] = 16'hffff;
  rom[09171] = 16'hffff;
  rom[09172] = 16'hffff;
  rom[09173] = 16'hffff;
  rom[09174] = 16'hffff;
  rom[09175] = 16'hffff;
  rom[09176] = 16'hffff;
  rom[09177] = 16'hffff;
  rom[09178] = 16'hffff;
  rom[09179] = 16'hffff;
  rom[09180] = 16'hffff;
  rom[09181] = 16'hffff;
  rom[09182] = 16'hffff;
  rom[09183] = 16'hffff;
  rom[09184] = 16'hffff;
  rom[09185] = 16'hffff;
  rom[09186] = 16'hffff;
  rom[09187] = 16'hffff;
  rom[09188] = 16'hffff;
  rom[09189] = 16'hffff;
  rom[09190] = 16'hffff;
  rom[09191] = 16'hffff;
  rom[09192] = 16'hffff;
  rom[09193] = 16'hffff;
  rom[09194] = 16'hffff;
  rom[09195] = 16'hffff;
  rom[09196] = 16'hffff;
  rom[09197] = 16'hffff;
  rom[09198] = 16'hffff;
  rom[09199] = 16'hffff;
  rom[09200] = 16'hffff;
  rom[09201] = 16'hffff;
  rom[09202] = 16'hffff;
  rom[09203] = 16'hffff;
  rom[09204] = 16'hffff;
  rom[09205] = 16'hffff;
  rom[09206] = 16'hffff;
  rom[09207] = 16'hffff;
  rom[09208] = 16'hffff;
  rom[09209] = 16'hffff;
  rom[09210] = 16'hffff;
  rom[09211] = 16'hffff;
  rom[09212] = 16'hffff;
  rom[09213] = 16'hffff;
  rom[09214] = 16'hffff;
  rom[09215] = 16'hffff;
  rom[09216] = 16'hffff;
  rom[09217] = 16'hffff;
  rom[09218] = 16'hffff;
  rom[09219] = 16'hffff;
  rom[09220] = 16'hffff;
  rom[09221] = 16'hffff;
  rom[09222] = 16'hffff;
  rom[09223] = 16'hffff;
  rom[09224] = 16'hffff;
  rom[09225] = 16'hffff;
  rom[09226] = 16'hffff;
  rom[09227] = 16'hffff;
  rom[09228] = 16'hffff;
  rom[09229] = 16'hffff;
  rom[09230] = 16'hffff;
  rom[09231] = 16'hffff;
  rom[09232] = 16'hffff;
  rom[09233] = 16'hffff;
  rom[09234] = 16'hffff;
  rom[09235] = 16'hffff;
  rom[09236] = 16'hffff;
  rom[09237] = 16'hffff;
  rom[09238] = 16'hffff;
  rom[09239] = 16'hffff;
  rom[09240] = 16'hffff;
  rom[09241] = 16'hffff;
  rom[09242] = 16'hffff;
  rom[09243] = 16'hffff;
  rom[09244] = 16'hffff;
  rom[09245] = 16'hffff;
  rom[09246] = 16'hffff;
  rom[09247] = 16'hff5c;
  rom[09248] = 16'h93aa;
  rom[09249] = 16'ha3e8;
  rom[09250] = 16'hdd8a;
  rom[09251] = 16'hed89;
  rom[09252] = 16'hfd48;
  rom[09253] = 16'hfd29;
  rom[09254] = 16'hf508;
  rom[09255] = 16'hfd69;
  rom[09256] = 16'hfd88;
  rom[09257] = 16'hfda7;
  rom[09258] = 16'hf567;
  rom[09259] = 16'hf58a;
  rom[09260] = 16'he58c;
  rom[09261] = 16'hb42a;
  rom[09262] = 16'h3921;
  rom[09263] = 16'h20a1;
  rom[09264] = 16'h18a2;
  rom[09265] = 16'h18c3;
  rom[09266] = 16'h1082;
  rom[09267] = 16'h18a2;
  rom[09268] = 16'h18a2;
  rom[09269] = 16'h18a3;
  rom[09270] = 16'h1083;
  rom[09271] = 16'h10a4;
  rom[09272] = 16'h18a3;
  rom[09273] = 16'h20a1;
  rom[09274] = 16'h51e2;
  rom[09275] = 16'hcd2b;
  rom[09276] = 16'hedeb;
  rom[09277] = 16'hf5c9;
  rom[09278] = 16'hf5c8;
  rom[09279] = 16'hfde8;
  rom[09280] = 16'hfde8;
  rom[09281] = 16'hfde9;
  rom[09282] = 16'hf5e9;
  rom[09283] = 16'hfde8;
  rom[09284] = 16'hfe09;
  rom[09285] = 16'hfe08;
  rom[09286] = 16'hf607;
  rom[09287] = 16'hfe29;
  rom[09288] = 16'hf629;
  rom[09289] = 16'hfe2a;
  rom[09290] = 16'hf609;
  rom[09291] = 16'hfe29;
  rom[09292] = 16'hf609;
  rom[09293] = 16'hfe2a;
  rom[09294] = 16'hf609;
  rom[09295] = 16'hfe29;
  rom[09296] = 16'hfe09;
  rom[09297] = 16'hfe29;
  rom[09298] = 16'hf608;
  rom[09299] = 16'hfe29;
  rom[09300] = 16'hfe0a;
  rom[09301] = 16'hfe2a;
  rom[09302] = 16'hf609;
  rom[09303] = 16'hfe09;
  rom[09304] = 16'hfe09;
  rom[09305] = 16'hf5e9;
  rom[09306] = 16'hfe09;
  rom[09307] = 16'hfe09;
  rom[09308] = 16'hfe08;
  rom[09309] = 16'hfe09;
  rom[09310] = 16'hf5e8;
  rom[09311] = 16'hfe08;
  rom[09312] = 16'hf5e9;
  rom[09313] = 16'hf609;
  rom[09314] = 16'hfe29;
  rom[09315] = 16'hf5e7;
  rom[09316] = 16'hf608;
  rom[09317] = 16'hf5eb;
  rom[09318] = 16'hbc8a;
  rom[09319] = 16'h4101;
  rom[09320] = 16'h2061;
  rom[09321] = 16'h1062;
  rom[09322] = 16'h18c3;
  rom[09323] = 16'h10c2;
  rom[09324] = 16'h10c3;
  rom[09325] = 16'h1082;
  rom[09326] = 16'h10a2;
  rom[09327] = 16'h18a2;
  rom[09328] = 16'h10a3;
  rom[09329] = 16'h18a3;
  rom[09330] = 16'h1882;
  rom[09331] = 16'h30e1;
  rom[09332] = 16'h9bc8;
  rom[09333] = 16'hed8b;
  rom[09334] = 16'hf5c8;
  rom[09335] = 16'hfd68;
  rom[09336] = 16'hfd49;
  rom[09337] = 16'hfd68;
  rom[09338] = 16'hf588;
  rom[09339] = 16'hfd68;
  rom[09340] = 16'hfd69;
  rom[09341] = 16'hfd69;
  rom[09342] = 16'hf547;
  rom[09343] = 16'hf587;
  rom[09344] = 16'hed68;
  rom[09345] = 16'he5ad;
  rom[09346] = 16'h72c5;
  rom[09347] = 16'hde78;
  rom[09348] = 16'hffdf;
  rom[09349] = 16'hffff;
  rom[09350] = 16'he71c;
  rom[09351] = 16'h7b6d;
  rom[09352] = 16'hd659;
  rom[09353] = 16'hffff;
  rom[09354] = 16'hffff;
  rom[09355] = 16'hffff;
  rom[09356] = 16'hffff;
  rom[09357] = 16'hffff;
  rom[09358] = 16'hffff;
  rom[09359] = 16'hffff;
  rom[09360] = 16'hffff;
  rom[09361] = 16'hffff;
  rom[09362] = 16'hffff;
  rom[09363] = 16'hffff;
  rom[09364] = 16'hffff;
  rom[09365] = 16'hffff;
  rom[09366] = 16'hffff;
  rom[09367] = 16'hffff;
  rom[09368] = 16'hffff;
  rom[09369] = 16'hffff;
  rom[09370] = 16'hffff;
  rom[09371] = 16'hffff;
  rom[09372] = 16'hffff;
  rom[09373] = 16'hffff;
  rom[09374] = 16'hffff;
  rom[09375] = 16'hffff;
  rom[09376] = 16'hffff;
  rom[09377] = 16'hffff;
  rom[09378] = 16'hffff;
  rom[09379] = 16'hffff;
  rom[09380] = 16'hffff;
  rom[09381] = 16'hffff;
  rom[09382] = 16'hffff;
  rom[09383] = 16'hffff;
  rom[09384] = 16'hffff;
  rom[09385] = 16'hffff;
  rom[09386] = 16'hffff;
  rom[09387] = 16'hffff;
  rom[09388] = 16'hffff;
  rom[09389] = 16'hffff;
  rom[09390] = 16'hffff;
  rom[09391] = 16'hffff;
  rom[09392] = 16'hffff;
  rom[09393] = 16'hffff;
  rom[09394] = 16'hffff;
  rom[09395] = 16'hffff;
  rom[09396] = 16'hffff;
  rom[09397] = 16'hffff;
  rom[09398] = 16'hffff;
  rom[09399] = 16'hffff;
  rom[09400] = 16'hffff;
  rom[09401] = 16'hffff;
  rom[09402] = 16'hffff;
  rom[09403] = 16'hffff;
  rom[09404] = 16'hffff;
  rom[09405] = 16'hffff;
  rom[09406] = 16'hffff;
  rom[09407] = 16'hffff;
  rom[09408] = 16'hffff;
  rom[09409] = 16'hffff;
  rom[09410] = 16'hffff;
  rom[09411] = 16'hffff;
  rom[09412] = 16'hffff;
  rom[09413] = 16'hffff;
  rom[09414] = 16'hffff;
  rom[09415] = 16'hffff;
  rom[09416] = 16'hffff;
  rom[09417] = 16'hffff;
  rom[09418] = 16'hffff;
  rom[09419] = 16'hffff;
  rom[09420] = 16'hffff;
  rom[09421] = 16'hffff;
  rom[09422] = 16'hffff;
  rom[09423] = 16'hffff;
  rom[09424] = 16'hffff;
  rom[09425] = 16'hffff;
  rom[09426] = 16'hffff;
  rom[09427] = 16'hffff;
  rom[09428] = 16'hffff;
  rom[09429] = 16'hffff;
  rom[09430] = 16'hffff;
  rom[09431] = 16'hffff;
  rom[09432] = 16'hffff;
  rom[09433] = 16'hffff;
  rom[09434] = 16'hffff;
  rom[09435] = 16'hffff;
  rom[09436] = 16'hffff;
  rom[09437] = 16'hffff;
  rom[09438] = 16'hffff;
  rom[09439] = 16'hffff;
  rom[09440] = 16'hffff;
  rom[09441] = 16'hffff;
  rom[09442] = 16'hffff;
  rom[09443] = 16'hffff;
  rom[09444] = 16'hffff;
  rom[09445] = 16'hffff;
  rom[09446] = 16'hffdf;
  rom[09447] = 16'hacd1;
  rom[09448] = 16'h8b48;
  rom[09449] = 16'hcd2b;
  rom[09450] = 16'hed8a;
  rom[09451] = 16'hed88;
  rom[09452] = 16'hfd89;
  rom[09453] = 16'hfd49;
  rom[09454] = 16'hfd6a;
  rom[09455] = 16'hfd69;
  rom[09456] = 16'hfd88;
  rom[09457] = 16'hfd87;
  rom[09458] = 16'hfda7;
  rom[09459] = 16'hf587;
  rom[09460] = 16'hf5aa;
  rom[09461] = 16'he58c;
  rom[09462] = 16'ha3a9;
  rom[09463] = 16'h30c1;
  rom[09464] = 16'h20a2;
  rom[09465] = 16'h18a3;
  rom[09466] = 16'h18a3;
  rom[09467] = 16'h18c3;
  rom[09468] = 16'h18c3;
  rom[09469] = 16'h0841;
  rom[09470] = 16'h18c3;
  rom[09471] = 16'h10c3;
  rom[09472] = 16'h18c3;
  rom[09473] = 16'h18a0;
  rom[09474] = 16'h3101;
  rom[09475] = 16'h8347;
  rom[09476] = 16'hee0f;
  rom[09477] = 16'hedeb;
  rom[09478] = 16'hf5c9;
  rom[09479] = 16'hfe29;
  rom[09480] = 16'hfe49;
  rom[09481] = 16'hfe2a;
  rom[09482] = 16'hf5c9;
  rom[09483] = 16'hf5ea;
  rom[09484] = 16'hfe4b;
  rom[09485] = 16'hfe09;
  rom[09486] = 16'hfe09;
  rom[09487] = 16'hfe08;
  rom[09488] = 16'hfe4a;
  rom[09489] = 16'hfe09;
  rom[09490] = 16'hfe09;
  rom[09491] = 16'hf62a;
  rom[09492] = 16'hfe09;
  rom[09493] = 16'hfe2a;
  rom[09494] = 16'hfe29;
  rom[09495] = 16'hfe28;
  rom[09496] = 16'hfe29;
  rom[09497] = 16'hfe28;
  rom[09498] = 16'hfe29;
  rom[09499] = 16'hfe28;
  rom[09500] = 16'hfe29;
  rom[09501] = 16'hfe09;
  rom[09502] = 16'hf62a;
  rom[09503] = 16'hfe08;
  rom[09504] = 16'hfe09;
  rom[09505] = 16'hfe28;
  rom[09506] = 16'hfe08;
  rom[09507] = 16'hfe08;
  rom[09508] = 16'hfe09;
  rom[09509] = 16'hf5e9;
  rom[09510] = 16'hfe2a;
  rom[09511] = 16'hfe0a;
  rom[09512] = 16'hedc9;
  rom[09513] = 16'hf60a;
  rom[09514] = 16'hf5e9;
  rom[09515] = 16'hf609;
  rom[09516] = 16'hf5ea;
  rom[09517] = 16'hedcd;
  rom[09518] = 16'h82e6;
  rom[09519] = 16'h2040;
  rom[09520] = 16'h28c4;
  rom[09521] = 16'h1083;
  rom[09522] = 16'h18e4;
  rom[09523] = 16'h10c2;
  rom[09524] = 16'h10c2;
  rom[09525] = 16'h10a2;
  rom[09526] = 16'h10c3;
  rom[09527] = 16'h10c3;
  rom[09528] = 16'h10a3;
  rom[09529] = 16'h18a3;
  rom[09530] = 16'h28c2;
  rom[09531] = 16'h93aa;
  rom[09532] = 16'hdd4c;
  rom[09533] = 16'hfdeb;
  rom[09534] = 16'hfd86;
  rom[09535] = 16'hfda8;
  rom[09536] = 16'hfd69;
  rom[09537] = 16'hfd89;
  rom[09538] = 16'hf569;
  rom[09539] = 16'hfd88;
  rom[09540] = 16'hfd69;
  rom[09541] = 16'hfd49;
  rom[09542] = 16'hfd68;
  rom[09543] = 16'hf587;
  rom[09544] = 16'hf5a9;
  rom[09545] = 16'he58c;
  rom[09546] = 16'hac0a;
  rom[09547] = 16'h9c2e;
  rom[09548] = 16'hffff;
  rom[09549] = 16'hffdf;
  rom[09550] = 16'hffbf;
  rom[09551] = 16'h83cf;
  rom[09552] = 16'h9c92;
  rom[09553] = 16'hffff;
  rom[09554] = 16'hffff;
  rom[09555] = 16'hffdf;
  rom[09556] = 16'hffff;
  rom[09557] = 16'hffdf;
  rom[09558] = 16'hffff;
  rom[09559] = 16'hffff;
  rom[09560] = 16'hffff;
  rom[09561] = 16'hffff;
  rom[09562] = 16'hffff;
  rom[09563] = 16'hffff;
  rom[09564] = 16'hffff;
  rom[09565] = 16'hffff;
  rom[09566] = 16'hffff;
  rom[09567] = 16'hffff;
  rom[09568] = 16'hffff;
  rom[09569] = 16'hffff;
  rom[09570] = 16'hffff;
  rom[09571] = 16'hffff;
  rom[09572] = 16'hffff;
  rom[09573] = 16'hffff;
  rom[09574] = 16'hffff;
  rom[09575] = 16'hffff;
  rom[09576] = 16'hffff;
  rom[09577] = 16'hffff;
  rom[09578] = 16'hffff;
  rom[09579] = 16'hffff;
  rom[09580] = 16'hffff;
  rom[09581] = 16'hffff;
  rom[09582] = 16'hffff;
  rom[09583] = 16'hffff;
  rom[09584] = 16'hffff;
  rom[09585] = 16'hffff;
  rom[09586] = 16'hffff;
  rom[09587] = 16'hffff;
  rom[09588] = 16'hffff;
  rom[09589] = 16'hffff;
  rom[09590] = 16'hffff;
  rom[09591] = 16'hffff;
  rom[09592] = 16'hffff;
  rom[09593] = 16'hffff;
  rom[09594] = 16'hffff;
  rom[09595] = 16'hffff;
  rom[09596] = 16'hffff;
  rom[09597] = 16'hffff;
  rom[09598] = 16'hffff;
  rom[09599] = 16'hffff;
  rom[09600] = 16'hffff;
  rom[09601] = 16'hffff;
  rom[09602] = 16'hffff;
  rom[09603] = 16'hffff;
  rom[09604] = 16'hffff;
  rom[09605] = 16'hffff;
  rom[09606] = 16'hffff;
  rom[09607] = 16'hffff;
  rom[09608] = 16'hffff;
  rom[09609] = 16'hffff;
  rom[09610] = 16'hffff;
  rom[09611] = 16'hffff;
  rom[09612] = 16'hffff;
  rom[09613] = 16'hffff;
  rom[09614] = 16'hffff;
  rom[09615] = 16'hffff;
  rom[09616] = 16'hffff;
  rom[09617] = 16'hffff;
  rom[09618] = 16'hffff;
  rom[09619] = 16'hffff;
  rom[09620] = 16'hffff;
  rom[09621] = 16'hffff;
  rom[09622] = 16'hffff;
  rom[09623] = 16'hffff;
  rom[09624] = 16'hffff;
  rom[09625] = 16'hffff;
  rom[09626] = 16'hffff;
  rom[09627] = 16'hffff;
  rom[09628] = 16'hffff;
  rom[09629] = 16'hffff;
  rom[09630] = 16'hffff;
  rom[09631] = 16'hffff;
  rom[09632] = 16'hffff;
  rom[09633] = 16'hffff;
  rom[09634] = 16'hffff;
  rom[09635] = 16'hffff;
  rom[09636] = 16'hffff;
  rom[09637] = 16'hffff;
  rom[09638] = 16'hffff;
  rom[09639] = 16'hffff;
  rom[09640] = 16'hffff;
  rom[09641] = 16'hffff;
  rom[09642] = 16'hffff;
  rom[09643] = 16'hffff;
  rom[09644] = 16'hffff;
  rom[09645] = 16'hffff;
  rom[09646] = 16'he6da;
  rom[09647] = 16'h8b8b;
  rom[09648] = 16'hac29;
  rom[09649] = 16'he5ab;
  rom[09650] = 16'hed88;
  rom[09651] = 16'hf588;
  rom[09652] = 16'hf528;
  rom[09653] = 16'hfd29;
  rom[09654] = 16'hfd28;
  rom[09655] = 16'hfd89;
  rom[09656] = 16'hf588;
  rom[09657] = 16'hfd87;
  rom[09658] = 16'hfda7;
  rom[09659] = 16'hfd66;
  rom[09660] = 16'hf587;
  rom[09661] = 16'hf5ab;
  rom[09662] = 16'hd50c;
  rom[09663] = 16'h7aa6;
  rom[09664] = 16'h2060;
  rom[09665] = 16'h20a2;
  rom[09666] = 16'h1882;
  rom[09667] = 16'h1062;
  rom[09668] = 16'h18a3;
  rom[09669] = 16'h10a2;
  rom[09670] = 16'h10c2;
  rom[09671] = 16'h1081;
  rom[09672] = 16'h10c1;
  rom[09673] = 16'h10a1;
  rom[09674] = 16'h1060;
  rom[09675] = 16'h51c3;
  rom[09676] = 16'hb4ed;
  rom[09677] = 16'he60e;
  rom[09678] = 16'hee2d;
  rom[09679] = 16'hedea;
  rom[09680] = 16'he5c9;
  rom[09681] = 16'hedeb;
  rom[09682] = 16'hfe6d;
  rom[09683] = 16'hf60c;
  rom[09684] = 16'hedca;
  rom[09685] = 16'hf62a;
  rom[09686] = 16'hfe4a;
  rom[09687] = 16'hfe09;
  rom[09688] = 16'hedc8;
  rom[09689] = 16'hfe4a;
  rom[09690] = 16'hfe49;
  rom[09691] = 16'hf5e8;
  rom[09692] = 16'hf629;
  rom[09693] = 16'hf608;
  rom[09694] = 16'hfe29;
  rom[09695] = 16'hfe29;
  rom[09696] = 16'hf609;
  rom[09697] = 16'hfe29;
  rom[09698] = 16'hfe08;
  rom[09699] = 16'hfe29;
  rom[09700] = 16'hf628;
  rom[09701] = 16'hfe29;
  rom[09702] = 16'hfe49;
  rom[09703] = 16'hfe49;
  rom[09704] = 16'hf628;
  rom[09705] = 16'hfe69;
  rom[09706] = 16'hf607;
  rom[09707] = 16'hf609;
  rom[09708] = 16'hfe29;
  rom[09709] = 16'hf60a;
  rom[09710] = 16'hedaa;
  rom[09711] = 16'hf5ec;
  rom[09712] = 16'hf62d;
  rom[09713] = 16'hedeb;
  rom[09714] = 16'hedeb;
  rom[09715] = 16'hf60d;
  rom[09716] = 16'hedee;
  rom[09717] = 16'hc4cc;
  rom[09718] = 16'h3901;
  rom[09719] = 16'h30e2;
  rom[09720] = 16'h1062;
  rom[09721] = 16'h1083;
  rom[09722] = 16'h10a3;
  rom[09723] = 16'h10e2;
  rom[09724] = 16'h10c2;
  rom[09725] = 16'h10c2;
  rom[09726] = 16'h0882;
  rom[09727] = 16'h10a3;
  rom[09728] = 16'h10c2;
  rom[09729] = 16'h18a0;
  rom[09730] = 16'h5a24;
  rom[09731] = 16'hd52e;
  rom[09732] = 16'hed8b;
  rom[09733] = 16'hfd89;
  rom[09734] = 16'hfd66;
  rom[09735] = 16'hfd88;
  rom[09736] = 16'hf547;
  rom[09737] = 16'hfda9;
  rom[09738] = 16'hf568;
  rom[09739] = 16'hfd89;
  rom[09740] = 16'hfd49;
  rom[09741] = 16'hfd69;
  rom[09742] = 16'hfd68;
  rom[09743] = 16'hf566;
  rom[09744] = 16'hf588;
  rom[09745] = 16'he52a;
  rom[09746] = 16'hd4ec;
  rom[09747] = 16'h82e7;
  rom[09748] = 16'heed9;
  rom[09749] = 16'hffff;
  rom[09750] = 16'hffbe;
  rom[09751] = 16'h9c91;
  rom[09752] = 16'h738e;
  rom[09753] = 16'hffbf;
  rom[09754] = 16'hffff;
  rom[09755] = 16'hffff;
  rom[09756] = 16'hffff;
  rom[09757] = 16'hffff;
  rom[09758] = 16'hffff;
  rom[09759] = 16'hffff;
  rom[09760] = 16'hffff;
  rom[09761] = 16'hffff;
  rom[09762] = 16'hffff;
  rom[09763] = 16'hffff;
  rom[09764] = 16'hffff;
  rom[09765] = 16'hffff;
  rom[09766] = 16'hffff;
  rom[09767] = 16'hffff;
  rom[09768] = 16'hffff;
  rom[09769] = 16'hffff;
  rom[09770] = 16'hffff;
  rom[09771] = 16'hffff;
  rom[09772] = 16'hffff;
  rom[09773] = 16'hffff;
  rom[09774] = 16'hffff;
  rom[09775] = 16'hffff;
  rom[09776] = 16'hffff;
  rom[09777] = 16'hffff;
  rom[09778] = 16'hffff;
  rom[09779] = 16'hffff;
  rom[09780] = 16'hffff;
  rom[09781] = 16'hffff;
  rom[09782] = 16'hffff;
  rom[09783] = 16'hffff;
  rom[09784] = 16'hffff;
  rom[09785] = 16'hffff;
  rom[09786] = 16'hffff;
  rom[09787] = 16'hffff;
  rom[09788] = 16'hffff;
  rom[09789] = 16'hffff;
  rom[09790] = 16'hffff;
  rom[09791] = 16'hffff;
  rom[09792] = 16'hffff;
  rom[09793] = 16'hffff;
  rom[09794] = 16'hffff;
  rom[09795] = 16'hffff;
  rom[09796] = 16'hffff;
  rom[09797] = 16'hffff;
  rom[09798] = 16'hffff;
  rom[09799] = 16'hffff;
  rom[09800] = 16'hffff;
  rom[09801] = 16'hffff;
  rom[09802] = 16'hffff;
  rom[09803] = 16'hffff;
  rom[09804] = 16'hffff;
  rom[09805] = 16'hffff;
  rom[09806] = 16'hffff;
  rom[09807] = 16'hffff;
  rom[09808] = 16'hffff;
  rom[09809] = 16'hffff;
  rom[09810] = 16'hffff;
  rom[09811] = 16'hffff;
  rom[09812] = 16'hffff;
  rom[09813] = 16'hffff;
  rom[09814] = 16'hffff;
  rom[09815] = 16'hffff;
  rom[09816] = 16'hffff;
  rom[09817] = 16'hffff;
  rom[09818] = 16'hffff;
  rom[09819] = 16'hffff;
  rom[09820] = 16'hffff;
  rom[09821] = 16'hffff;
  rom[09822] = 16'hffff;
  rom[09823] = 16'hffff;
  rom[09824] = 16'hffff;
  rom[09825] = 16'hffff;
  rom[09826] = 16'hffff;
  rom[09827] = 16'hffff;
  rom[09828] = 16'hffff;
  rom[09829] = 16'hffff;
  rom[09830] = 16'hffff;
  rom[09831] = 16'hffff;
  rom[09832] = 16'hffff;
  rom[09833] = 16'hffff;
  rom[09834] = 16'hffff;
  rom[09835] = 16'hffff;
  rom[09836] = 16'hffff;
  rom[09837] = 16'hffff;
  rom[09838] = 16'hffff;
  rom[09839] = 16'hffff;
  rom[09840] = 16'hffff;
  rom[09841] = 16'hffff;
  rom[09842] = 16'hffff;
  rom[09843] = 16'hffff;
  rom[09844] = 16'hffff;
  rom[09845] = 16'hffff;
  rom[09846] = 16'hb4f2;
  rom[09847] = 16'h9ba9;
  rom[09848] = 16'hdd6c;
  rom[09849] = 16'he569;
  rom[09850] = 16'hfda8;
  rom[09851] = 16'hfd88;
  rom[09852] = 16'hfd48;
  rom[09853] = 16'hfd49;
  rom[09854] = 16'hfd6a;
  rom[09855] = 16'hf569;
  rom[09856] = 16'hfdaa;
  rom[09857] = 16'hf569;
  rom[09858] = 16'hfd89;
  rom[09859] = 16'hfd88;
  rom[09860] = 16'hfda9;
  rom[09861] = 16'hf569;
  rom[09862] = 16'hfdcd;
  rom[09863] = 16'hc4cb;
  rom[09864] = 16'h6a65;
  rom[09865] = 16'h1880;
  rom[09866] = 16'h18c2;
  rom[09867] = 16'h1082;
  rom[09868] = 16'h18a4;
  rom[09869] = 16'h18c3;
  rom[09870] = 16'h18e3;
  rom[09871] = 16'h08a1;
  rom[09872] = 16'h18e2;
  rom[09873] = 16'h10c2;
  rom[09874] = 16'h1882;
  rom[09875] = 16'h20c1;
  rom[09876] = 16'h7308;
  rom[09877] = 16'hac8b;
  rom[09878] = 16'hb48a;
  rom[09879] = 16'hbca9;
  rom[09880] = 16'hc4ea;
  rom[09881] = 16'hcd2b;
  rom[09882] = 16'hd58c;
  rom[09883] = 16'hddcd;
  rom[09884] = 16'hee0e;
  rom[09885] = 16'he60c;
  rom[09886] = 16'hedec;
  rom[09887] = 16'hf64b;
  rom[09888] = 16'hf62a;
  rom[09889] = 16'hf629;
  rom[09890] = 16'hfe6a;
  rom[09891] = 16'hf649;
  rom[09892] = 16'hfe49;
  rom[09893] = 16'hfe28;
  rom[09894] = 16'hfe29;
  rom[09895] = 16'hfe2a;
  rom[09896] = 16'hfe2a;
  rom[09897] = 16'hfe2a;
  rom[09898] = 16'hfe2a;
  rom[09899] = 16'hfe29;
  rom[09900] = 16'hfe49;
  rom[09901] = 16'hfe49;
  rom[09902] = 16'hfe29;
  rom[09903] = 16'hf629;
  rom[09904] = 16'hf649;
  rom[09905] = 16'hee29;
  rom[09906] = 16'hfe4b;
  rom[09907] = 16'hf62b;
  rom[09908] = 16'hf62c;
  rom[09909] = 16'hee2d;
  rom[09910] = 16'hedee;
  rom[09911] = 16'hd56c;
  rom[09912] = 16'hd56c;
  rom[09913] = 16'hcd0a;
  rom[09914] = 16'hbcaa;
  rom[09915] = 16'hb449;
  rom[09916] = 16'hb46c;
  rom[09917] = 16'h6a86;
  rom[09918] = 16'h28c1;
  rom[09919] = 16'h18c2;
  rom[09920] = 16'h10a2;
  rom[09921] = 16'h10c3;
  rom[09922] = 16'h18c4;
  rom[09923] = 16'h10c2;
  rom[09924] = 16'h18c2;
  rom[09925] = 16'h10a1;
  rom[09926] = 16'h18a2;
  rom[09927] = 16'h18a2;
  rom[09928] = 16'h18a1;
  rom[09929] = 16'h5a23;
  rom[09930] = 16'hc4eb;
  rom[09931] = 16'hedab;
  rom[09932] = 16'hfdaa;
  rom[09933] = 16'hf568;
  rom[09934] = 16'hfd89;
  rom[09935] = 16'hfda9;
  rom[09936] = 16'hfd88;
  rom[09937] = 16'hf588;
  rom[09938] = 16'hfda9;
  rom[09939] = 16'hf568;
  rom[09940] = 16'hfd89;
  rom[09941] = 16'hfd49;
  rom[09942] = 16'hfd89;
  rom[09943] = 16'hece5;
  rom[09944] = 16'hfda9;
  rom[09945] = 16'hed49;
  rom[09946] = 16'hed6d;
  rom[09947] = 16'h9b47;
  rom[09948] = 16'hac8f;
  rom[09949] = 16'hffdd;
  rom[09950] = 16'hffff;
  rom[09951] = 16'had35;
  rom[09952] = 16'h5acb;
  rom[09953] = 16'hd69a;
  rom[09954] = 16'hffff;
  rom[09955] = 16'hffff;
  rom[09956] = 16'hffff;
  rom[09957] = 16'hffff;
  rom[09958] = 16'hffff;
  rom[09959] = 16'hffff;
  rom[09960] = 16'hffff;
  rom[09961] = 16'hffff;
  rom[09962] = 16'hffff;
  rom[09963] = 16'hffff;
  rom[09964] = 16'hffff;
  rom[09965] = 16'hffff;
  rom[09966] = 16'hffff;
  rom[09967] = 16'hffff;
  rom[09968] = 16'hffff;
  rom[09969] = 16'hffff;
  rom[09970] = 16'hffff;
  rom[09971] = 16'hffff;
  rom[09972] = 16'hffff;
  rom[09973] = 16'hffff;
  rom[09974] = 16'hffff;
  rom[09975] = 16'hffff;
  rom[09976] = 16'hffff;
  rom[09977] = 16'hffff;
  rom[09978] = 16'hffff;
  rom[09979] = 16'hffff;
  rom[09980] = 16'hffff;
  rom[09981] = 16'hffff;
  rom[09982] = 16'hffff;
  rom[09983] = 16'hffff;
  rom[09984] = 16'hffff;
  rom[09985] = 16'hffff;
  rom[09986] = 16'hffff;
  rom[09987] = 16'hffff;
  rom[09988] = 16'hffff;
  rom[09989] = 16'hffff;
  rom[09990] = 16'hffff;
  rom[09991] = 16'hffff;
  rom[09992] = 16'hffff;
  rom[09993] = 16'hffff;
  rom[09994] = 16'hffff;
  rom[09995] = 16'hffff;
  rom[09996] = 16'hffff;
  rom[09997] = 16'hffff;
  rom[09998] = 16'hffff;
  rom[09999] = 16'hffff;
  rom[10000] = 16'hffff;
  rom[10001] = 16'hffff;
  rom[10002] = 16'hffff;
  rom[10003] = 16'hffff;
  rom[10004] = 16'hffff;
  rom[10005] = 16'hffff;
  rom[10006] = 16'hffff;
  rom[10007] = 16'hffff;
  rom[10008] = 16'hffff;
  rom[10009] = 16'hffff;
  rom[10010] = 16'hffff;
  rom[10011] = 16'hffff;
  rom[10012] = 16'hffff;
  rom[10013] = 16'hffff;
  rom[10014] = 16'hffff;
  rom[10015] = 16'hffff;
  rom[10016] = 16'hffff;
  rom[10017] = 16'hffff;
  rom[10018] = 16'hffff;
  rom[10019] = 16'hffff;
  rom[10020] = 16'hffff;
  rom[10021] = 16'hffff;
  rom[10022] = 16'hffff;
  rom[10023] = 16'hffff;
  rom[10024] = 16'hffff;
  rom[10025] = 16'hffff;
  rom[10026] = 16'hffff;
  rom[10027] = 16'hffff;
  rom[10028] = 16'hffff;
  rom[10029] = 16'hffff;
  rom[10030] = 16'hffff;
  rom[10031] = 16'hffff;
  rom[10032] = 16'hffff;
  rom[10033] = 16'hffff;
  rom[10034] = 16'hffff;
  rom[10035] = 16'hffff;
  rom[10036] = 16'hffff;
  rom[10037] = 16'hffff;
  rom[10038] = 16'hffff;
  rom[10039] = 16'hffff;
  rom[10040] = 16'hffff;
  rom[10041] = 16'hffff;
  rom[10042] = 16'hffff;
  rom[10043] = 16'hffff;
  rom[10044] = 16'hffff;
  rom[10045] = 16'hf71b;
  rom[10046] = 16'h8329;
  rom[10047] = 16'hc48c;
  rom[10048] = 16'hed8c;
  rom[10049] = 16'hf589;
  rom[10050] = 16'hf587;
  rom[10051] = 16'hfd68;
  rom[10052] = 16'hfd48;
  rom[10053] = 16'hfd49;
  rom[10054] = 16'hfd69;
  rom[10055] = 16'hfda9;
  rom[10056] = 16'hf588;
  rom[10057] = 16'hfdca;
  rom[10058] = 16'hed48;
  rom[10059] = 16'hfd8a;
  rom[10060] = 16'hfd89;
  rom[10061] = 16'hfd89;
  rom[10062] = 16'hed89;
  rom[10063] = 16'hee0c;
  rom[10064] = 16'hbcca;
  rom[10065] = 16'h5203;
  rom[10066] = 16'h1060;
  rom[10067] = 16'h2105;
  rom[10068] = 16'h18a3;
  rom[10069] = 16'h18c3;
  rom[10070] = 16'h0881;
  rom[10071] = 16'h10a2;
  rom[10072] = 16'h10e3;
  rom[10073] = 16'h18e4;
  rom[10074] = 16'h39c8;
  rom[10075] = 16'h6b0c;
  rom[10076] = 16'h734b;
  rom[10077] = 16'h8bec;
  rom[10078] = 16'h83c9;
  rom[10079] = 16'h93aa;
  rom[10080] = 16'h93c9;
  rom[10081] = 16'h93a9;
  rom[10082] = 16'h8347;
  rom[10083] = 16'h6263;
  rom[10084] = 16'h7b25;
  rom[10085] = 16'hac69;
  rom[10086] = 16'hddcd;
  rom[10087] = 16'hee4e;
  rom[10088] = 16'hf60c;
  rom[10089] = 16'hf62b;
  rom[10090] = 16'hf64b;
  rom[10091] = 16'hf66a;
  rom[10092] = 16'hf629;
  rom[10093] = 16'hfe69;
  rom[10094] = 16'hf609;
  rom[10095] = 16'hfe29;
  rom[10096] = 16'hfe0a;
  rom[10097] = 16'hfe2a;
  rom[10098] = 16'hf60a;
  rom[10099] = 16'hfe2a;
  rom[10100] = 16'hfe29;
  rom[10101] = 16'hfe29;
  rom[10102] = 16'hf62a;
  rom[10103] = 16'hfe6a;
  rom[10104] = 16'hf62b;
  rom[10105] = 16'hf64c;
  rom[10106] = 16'he60c;
  rom[10107] = 16'he5ed;
  rom[10108] = 16'hbcca;
  rom[10109] = 16'h93a7;
  rom[10110] = 16'h72a3;
  rom[10111] = 16'h7ae5;
  rom[10112] = 16'h8b88;
  rom[10113] = 16'h93a9;
  rom[10114] = 16'h93c9;
  rom[10115] = 16'h93cb;
  rom[10116] = 16'h8bab;
  rom[10117] = 16'h7b4b;
  rom[10118] = 16'h736d;
  rom[10119] = 16'h52a9;
  rom[10120] = 16'h3186;
  rom[10121] = 16'h1904;
  rom[10122] = 16'h18e3;
  rom[10123] = 16'h10a2;
  rom[10124] = 16'h1041;
  rom[10125] = 16'h2904;
  rom[10126] = 16'h18a2;
  rom[10127] = 16'h1060;
  rom[10128] = 16'h49e3;
  rom[10129] = 16'hbcaa;
  rom[10130] = 16'he5aa;
  rom[10131] = 16'hf5c8;
  rom[10132] = 16'hf587;
  rom[10133] = 16'hfd88;
  rom[10134] = 16'hed69;
  rom[10135] = 16'hf589;
  rom[10136] = 16'hfdc9;
  rom[10137] = 16'hf587;
  rom[10138] = 16'hf588;
  rom[10139] = 16'hfd89;
  rom[10140] = 16'hfd49;
  rom[10141] = 16'hfd69;
  rom[10142] = 16'hf527;
  rom[10143] = 16'hfdc8;
  rom[10144] = 16'hf547;
  rom[10145] = 16'hfdaa;
  rom[10146] = 16'hdce9;
  rom[10147] = 16'hd4cc;
  rom[10148] = 16'h7ae7;
  rom[10149] = 16'hef1a;
  rom[10150] = 16'hffff;
  rom[10151] = 16'hb596;
  rom[10152] = 16'h2925;
  rom[10153] = 16'hbdb7;
  rom[10154] = 16'hffff;
  rom[10155] = 16'hffff;
  rom[10156] = 16'hffff;
  rom[10157] = 16'hffff;
  rom[10158] = 16'hffff;
  rom[10159] = 16'hffff;
  rom[10160] = 16'hffff;
  rom[10161] = 16'hffff;
  rom[10162] = 16'hffff;
  rom[10163] = 16'hffff;
  rom[10164] = 16'hffff;
  rom[10165] = 16'hffff;
  rom[10166] = 16'hffff;
  rom[10167] = 16'hffff;
  rom[10168] = 16'hffff;
  rom[10169] = 16'hffff;
  rom[10170] = 16'hffff;
  rom[10171] = 16'hffff;
  rom[10172] = 16'hffff;
  rom[10173] = 16'hffff;
  rom[10174] = 16'hffff;
  rom[10175] = 16'hffff;
  rom[10176] = 16'hffff;
  rom[10177] = 16'hffff;
  rom[10178] = 16'hffff;
  rom[10179] = 16'hffff;
  rom[10180] = 16'hffff;
  rom[10181] = 16'hffff;
  rom[10182] = 16'hffff;
  rom[10183] = 16'hffff;
  rom[10184] = 16'hffff;
  rom[10185] = 16'hffff;
  rom[10186] = 16'hffff;
  rom[10187] = 16'hffff;
  rom[10188] = 16'hffff;
  rom[10189] = 16'hffff;
  rom[10190] = 16'hffff;
  rom[10191] = 16'hffff;
  rom[10192] = 16'hffff;
  rom[10193] = 16'hffff;
  rom[10194] = 16'hffff;
  rom[10195] = 16'hffff;
  rom[10196] = 16'hffff;
  rom[10197] = 16'hffff;
  rom[10198] = 16'hffff;
  rom[10199] = 16'hffff;
  rom[10200] = 16'hffff;
  rom[10201] = 16'hffff;
  rom[10202] = 16'hffff;
  rom[10203] = 16'hffff;
  rom[10204] = 16'hffff;
  rom[10205] = 16'hffff;
  rom[10206] = 16'hffff;
  rom[10207] = 16'hffff;
  rom[10208] = 16'hffff;
  rom[10209] = 16'hffff;
  rom[10210] = 16'hffff;
  rom[10211] = 16'hffff;
  rom[10212] = 16'hffff;
  rom[10213] = 16'hffff;
  rom[10214] = 16'hffff;
  rom[10215] = 16'hffff;
  rom[10216] = 16'hffff;
  rom[10217] = 16'hffff;
  rom[10218] = 16'hffff;
  rom[10219] = 16'hffff;
  rom[10220] = 16'hffff;
  rom[10221] = 16'hffff;
  rom[10222] = 16'hffff;
  rom[10223] = 16'hffff;
  rom[10224] = 16'hffff;
  rom[10225] = 16'hffff;
  rom[10226] = 16'hffff;
  rom[10227] = 16'hffff;
  rom[10228] = 16'hffff;
  rom[10229] = 16'hffff;
  rom[10230] = 16'hffff;
  rom[10231] = 16'hffff;
  rom[10232] = 16'hffff;
  rom[10233] = 16'hffff;
  rom[10234] = 16'hffff;
  rom[10235] = 16'hffff;
  rom[10236] = 16'hffff;
  rom[10237] = 16'hffff;
  rom[10238] = 16'hffff;
  rom[10239] = 16'hffff;
  rom[10240] = 16'hffff;
  rom[10241] = 16'hffff;
  rom[10242] = 16'hffff;
  rom[10243] = 16'hffdf;
  rom[10244] = 16'hffbe;
  rom[10245] = 16'hb4f2;
  rom[10246] = 16'h9349;
  rom[10247] = 16'hdd0c;
  rom[10248] = 16'hf56a;
  rom[10249] = 16'hfd88;
  rom[10250] = 16'hfd66;
  rom[10251] = 16'hfd67;
  rom[10252] = 16'hfd49;
  rom[10253] = 16'hfd49;
  rom[10254] = 16'hfd6a;
  rom[10255] = 16'hfd89;
  rom[10256] = 16'hfdaa;
  rom[10257] = 16'hed68;
  rom[10258] = 16'hfdaa;
  rom[10259] = 16'hf569;
  rom[10260] = 16'hfd8a;
  rom[10261] = 16'hfd89;
  rom[10262] = 16'hfdc9;
  rom[10263] = 16'hed89;
  rom[10264] = 16'hee2e;
  rom[10265] = 16'hacac;
  rom[10266] = 16'h49e5;
  rom[10267] = 16'h1061;
  rom[10268] = 16'h18c3;
  rom[10269] = 16'h2965;
  rom[10270] = 16'h52aa;
  rom[10271] = 16'h7c10;
  rom[10272] = 16'had56;
  rom[10273] = 16'hbdf8;
  rom[10274] = 16'he71d;
  rom[10275] = 16'hef3d;
  rom[10276] = 16'hf75d;
  rom[10277] = 16'hf79c;
  rom[10278] = 16'hffbd;
  rom[10279] = 16'hffbd;
  rom[10280] = 16'hff5b;
  rom[10281] = 16'hef1a;
  rom[10282] = 16'heefa;
  rom[10283] = 16'hd656;
  rom[10284] = 16'hc593;
  rom[10285] = 16'ha4ae;
  rom[10286] = 16'h8b88;
  rom[10287] = 16'h8ba7;
  rom[10288] = 16'hac89;
  rom[10289] = 16'hd58c;
  rom[10290] = 16'he60d;
  rom[10291] = 16'hf66d;
  rom[10292] = 16'hf64b;
  rom[10293] = 16'hf64a;
  rom[10294] = 16'hfe4a;
  rom[10295] = 16'hfe29;
  rom[10296] = 16'hfe4a;
  rom[10297] = 16'hfe2a;
  rom[10298] = 16'hfe4a;
  rom[10299] = 16'hf629;
  rom[10300] = 16'hfe6b;
  rom[10301] = 16'hf62a;
  rom[10302] = 16'hf64c;
  rom[10303] = 16'hf64d;
  rom[10304] = 16'hddcc;
  rom[10305] = 16'hc50b;
  rom[10306] = 16'ha409;
  rom[10307] = 16'h8b67;
  rom[10308] = 16'h9c0b;
  rom[10309] = 16'hacef;
  rom[10310] = 16'hcdd4;
  rom[10311] = 16'hde76;
  rom[10312] = 16'hf75a;
  rom[10313] = 16'hf75a;
  rom[10314] = 16'hffdd;
  rom[10315] = 16'hff7c;
  rom[10316] = 16'hffbe;
  rom[10317] = 16'hf77c;
  rom[10318] = 16'hef5d;
  rom[10319] = 16'hdf3b;
  rom[10320] = 16'hd6da;
  rom[10321] = 16'had96;
  rom[10322] = 16'h94d3;
  rom[10323] = 16'h634d;
  rom[10324] = 16'h41e8;
  rom[10325] = 16'h2104;
  rom[10326] = 16'h1882;
  rom[10327] = 16'h49a5;
  rom[10328] = 16'hac8d;
  rom[10329] = 16'hddad;
  rom[10330] = 16'hf5ca;
  rom[10331] = 16'hfda7;
  rom[10332] = 16'hfdc7;
  rom[10333] = 16'hfdc9;
  rom[10334] = 16'hfd8a;
  rom[10335] = 16'hf589;
  rom[10336] = 16'hfda9;
  rom[10337] = 16'hfd88;
  rom[10338] = 16'hfd89;
  rom[10339] = 16'hf548;
  rom[10340] = 16'hfd6a;
  rom[10341] = 16'hfd68;
  rom[10342] = 16'hfd47;
  rom[10343] = 16'hfdc9;
  rom[10344] = 16'hf547;
  rom[10345] = 16'hfd88;
  rom[10346] = 16'hf56b;
  rom[10347] = 16'hdcec;
  rom[10348] = 16'h8b28;
  rom[10349] = 16'hc5d5;
  rom[10350] = 16'hffff;
  rom[10351] = 16'hbdf8;
  rom[10352] = 16'h2945;
  rom[10353] = 16'h9cb2;
  rom[10354] = 16'hffbe;
  rom[10355] = 16'hffff;
  rom[10356] = 16'hffff;
  rom[10357] = 16'hffff;
  rom[10358] = 16'hffff;
  rom[10359] = 16'hffff;
  rom[10360] = 16'hffff;
  rom[10361] = 16'hffff;
  rom[10362] = 16'hffff;
  rom[10363] = 16'hffff;
  rom[10364] = 16'hffff;
  rom[10365] = 16'hffff;
  rom[10366] = 16'hffff;
  rom[10367] = 16'hffff;
  rom[10368] = 16'hffff;
  rom[10369] = 16'hffff;
  rom[10370] = 16'hffff;
  rom[10371] = 16'hffff;
  rom[10372] = 16'hffff;
  rom[10373] = 16'hffff;
  rom[10374] = 16'hffff;
  rom[10375] = 16'hffff;
  rom[10376] = 16'hffff;
  rom[10377] = 16'hffff;
  rom[10378] = 16'hffff;
  rom[10379] = 16'hffff;
  rom[10380] = 16'hffff;
  rom[10381] = 16'hffff;
  rom[10382] = 16'hffff;
  rom[10383] = 16'hffff;
  rom[10384] = 16'hffff;
  rom[10385] = 16'hffff;
  rom[10386] = 16'hffff;
  rom[10387] = 16'hffff;
  rom[10388] = 16'hffff;
  rom[10389] = 16'hffff;
  rom[10390] = 16'hffff;
  rom[10391] = 16'hffff;
  rom[10392] = 16'hffff;
  rom[10393] = 16'hffff;
  rom[10394] = 16'hffff;
  rom[10395] = 16'hffff;
  rom[10396] = 16'hffff;
  rom[10397] = 16'hffff;
  rom[10398] = 16'hffff;
  rom[10399] = 16'hffff;
  rom[10400] = 16'hffff;
  rom[10401] = 16'hffff;
  rom[10402] = 16'hffff;
  rom[10403] = 16'hffff;
  rom[10404] = 16'hffff;
  rom[10405] = 16'hffff;
  rom[10406] = 16'hffff;
  rom[10407] = 16'hffff;
  rom[10408] = 16'hffff;
  rom[10409] = 16'hffff;
  rom[10410] = 16'hffff;
  rom[10411] = 16'hffff;
  rom[10412] = 16'hffff;
  rom[10413] = 16'hffff;
  rom[10414] = 16'hffff;
  rom[10415] = 16'hffff;
  rom[10416] = 16'hffff;
  rom[10417] = 16'hffff;
  rom[10418] = 16'hffff;
  rom[10419] = 16'hffff;
  rom[10420] = 16'hffff;
  rom[10421] = 16'hffff;
  rom[10422] = 16'hffff;
  rom[10423] = 16'hffff;
  rom[10424] = 16'hffff;
  rom[10425] = 16'hffff;
  rom[10426] = 16'hffff;
  rom[10427] = 16'hffff;
  rom[10428] = 16'hffff;
  rom[10429] = 16'hffff;
  rom[10430] = 16'hffff;
  rom[10431] = 16'hffff;
  rom[10432] = 16'hffff;
  rom[10433] = 16'hffff;
  rom[10434] = 16'hffff;
  rom[10435] = 16'hffff;
  rom[10436] = 16'hffff;
  rom[10437] = 16'hffff;
  rom[10438] = 16'hffff;
  rom[10439] = 16'hffff;
  rom[10440] = 16'hffff;
  rom[10441] = 16'hffff;
  rom[10442] = 16'hffdf;
  rom[10443] = 16'hffde;
  rom[10444] = 16'hef1a;
  rom[10445] = 16'h8b4a;
  rom[10446] = 16'hb42b;
  rom[10447] = 16'hf56d;
  rom[10448] = 16'hf528;
  rom[10449] = 16'hfd88;
  rom[10450] = 16'hf506;
  rom[10451] = 16'hfd89;
  rom[10452] = 16'hf549;
  rom[10453] = 16'hfd49;
  rom[10454] = 16'hfd49;
  rom[10455] = 16'hfd89;
  rom[10456] = 16'hf588;
  rom[10457] = 16'hfda8;
  rom[10458] = 16'hf587;
  rom[10459] = 16'hfdc9;
  rom[10460] = 16'hf567;
  rom[10461] = 16'hfda9;
  rom[10462] = 16'hf568;
  rom[10463] = 16'hfdec;
  rom[10464] = 16'hd54b;
  rom[10465] = 16'hcd4f;
  rom[10466] = 16'h6267;
  rom[10467] = 16'h3964;
  rom[10468] = 16'h7bcf;
  rom[10469] = 16'hc5f8;
  rom[10470] = 16'he73d;
  rom[10471] = 16'hf79f;
  rom[10472] = 16'hffdf;
  rom[10473] = 16'hffff;
  rom[10474] = 16'hffdf;
  rom[10475] = 16'hffdf;
  rom[10476] = 16'hffff;
  rom[10477] = 16'hffff;
  rom[10478] = 16'hffdf;
  rom[10479] = 16'hffff;
  rom[10480] = 16'hffff;
  rom[10481] = 16'hffff;
  rom[10482] = 16'hffff;
  rom[10483] = 16'hffff;
  rom[10484] = 16'hffde;
  rom[10485] = 16'hffbd;
  rom[10486] = 16'hf73b;
  rom[10487] = 16'hd615;
  rom[10488] = 16'h9c4d;
  rom[10489] = 16'h7b27;
  rom[10490] = 16'h93c8;
  rom[10491] = 16'hd5cf;
  rom[10492] = 16'he60d;
  rom[10493] = 16'hf66d;
  rom[10494] = 16'hf66a;
  rom[10495] = 16'hfe48;
  rom[10496] = 16'hfe67;
  rom[10497] = 16'hfe68;
  rom[10498] = 16'hf628;
  rom[10499] = 16'hf64a;
  rom[10500] = 16'hee4b;
  rom[10501] = 16'hee4d;
  rom[10502] = 16'hee4e;
  rom[10503] = 16'hbcea;
  rom[10504] = 16'h72e4;
  rom[10505] = 16'h8347;
  rom[10506] = 16'hc551;
  rom[10507] = 16'hf6f9;
  rom[10508] = 16'hf75c;
  rom[10509] = 16'hffde;
  rom[10510] = 16'hffdd;
  rom[10511] = 16'hffff;
  rom[10512] = 16'hfffe;
  rom[10513] = 16'hffff;
  rom[10514] = 16'hffff;
  rom[10515] = 16'hffff;
  rom[10516] = 16'hffff;
  rom[10517] = 16'hffff;
  rom[10518] = 16'hffff;
  rom[10519] = 16'hffff;
  rom[10520] = 16'hffff;
  rom[10521] = 16'hffff;
  rom[10522] = 16'hffdf;
  rom[10523] = 16'hf77f;
  rom[10524] = 16'hce9b;
  rom[10525] = 16'ha515;
  rom[10526] = 16'h524a;
  rom[10527] = 16'h5207;
  rom[10528] = 16'hb4ae;
  rom[10529] = 16'he5cf;
  rom[10530] = 16'he58a;
  rom[10531] = 16'hfdc8;
  rom[10532] = 16'hfda7;
  rom[10533] = 16'hf587;
  rom[10534] = 16'hf5a8;
  rom[10535] = 16'hf588;
  rom[10536] = 16'hf588;
  rom[10537] = 16'hf587;
  rom[10538] = 16'hfd89;
  rom[10539] = 16'hfd89;
  rom[10540] = 16'hfd48;
  rom[10541] = 16'hfd68;
  rom[10542] = 16'hf527;
  rom[10543] = 16'hfda9;
  rom[10544] = 16'hfd68;
  rom[10545] = 16'hf548;
  rom[10546] = 16'hf549;
  rom[10547] = 16'hf58d;
  rom[10548] = 16'hac2a;
  rom[10549] = 16'ha48f;
  rom[10550] = 16'hffbf;
  rom[10551] = 16'hce59;
  rom[10552] = 16'h4207;
  rom[10553] = 16'h8bae;
  rom[10554] = 16'hf77d;
  rom[10555] = 16'hffff;
  rom[10556] = 16'hffff;
  rom[10557] = 16'hffff;
  rom[10558] = 16'hffff;
  rom[10559] = 16'hffff;
  rom[10560] = 16'hffff;
  rom[10561] = 16'hffff;
  rom[10562] = 16'hffff;
  rom[10563] = 16'hffff;
  rom[10564] = 16'hffff;
  rom[10565] = 16'hffff;
  rom[10566] = 16'hffff;
  rom[10567] = 16'hffff;
  rom[10568] = 16'hffff;
  rom[10569] = 16'hffff;
  rom[10570] = 16'hffff;
  rom[10571] = 16'hffff;
  rom[10572] = 16'hffff;
  rom[10573] = 16'hffff;
  rom[10574] = 16'hffff;
  rom[10575] = 16'hffff;
  rom[10576] = 16'hffff;
  rom[10577] = 16'hffff;
  rom[10578] = 16'hffff;
  rom[10579] = 16'hffff;
  rom[10580] = 16'hffff;
  rom[10581] = 16'hffff;
  rom[10582] = 16'hffff;
  rom[10583] = 16'hffff;
  rom[10584] = 16'hffff;
  rom[10585] = 16'hffff;
  rom[10586] = 16'hffff;
  rom[10587] = 16'hffff;
  rom[10588] = 16'hffff;
  rom[10589] = 16'hffff;
  rom[10590] = 16'hffff;
  rom[10591] = 16'hffff;
  rom[10592] = 16'hffff;
  rom[10593] = 16'hffff;
  rom[10594] = 16'hffff;
  rom[10595] = 16'hffff;
  rom[10596] = 16'hffff;
  rom[10597] = 16'hffff;
  rom[10598] = 16'hffff;
  rom[10599] = 16'hffff;
  rom[10600] = 16'hffff;
  rom[10601] = 16'hffff;
  rom[10602] = 16'hffff;
  rom[10603] = 16'hffff;
  rom[10604] = 16'hffff;
  rom[10605] = 16'hffff;
  rom[10606] = 16'hffff;
  rom[10607] = 16'hffff;
  rom[10608] = 16'hffff;
  rom[10609] = 16'hffff;
  rom[10610] = 16'hffff;
  rom[10611] = 16'hffff;
  rom[10612] = 16'hffff;
  rom[10613] = 16'hffff;
  rom[10614] = 16'hffff;
  rom[10615] = 16'hffff;
  rom[10616] = 16'hffff;
  rom[10617] = 16'hffff;
  rom[10618] = 16'hffff;
  rom[10619] = 16'hffff;
  rom[10620] = 16'hffff;
  rom[10621] = 16'hffff;
  rom[10622] = 16'hffff;
  rom[10623] = 16'hffff;
  rom[10624] = 16'hffff;
  rom[10625] = 16'hffff;
  rom[10626] = 16'hffff;
  rom[10627] = 16'hffff;
  rom[10628] = 16'hffff;
  rom[10629] = 16'hffff;
  rom[10630] = 16'hffff;
  rom[10631] = 16'hffff;
  rom[10632] = 16'hffff;
  rom[10633] = 16'hffff;
  rom[10634] = 16'hffff;
  rom[10635] = 16'hffff;
  rom[10636] = 16'hffff;
  rom[10637] = 16'hffff;
  rom[10638] = 16'hffff;
  rom[10639] = 16'hffff;
  rom[10640] = 16'hffff;
  rom[10641] = 16'hffff;
  rom[10642] = 16'hffff;
  rom[10643] = 16'hfffe;
  rom[10644] = 16'hcdf5;
  rom[10645] = 16'h8b27;
  rom[10646] = 16'hdcec;
  rom[10647] = 16'hf56b;
  rom[10648] = 16'hfd68;
  rom[10649] = 16'hfd67;
  rom[10650] = 16'hfd48;
  rom[10651] = 16'hfd68;
  rom[10652] = 16'hfd69;
  rom[10653] = 16'hfd69;
  rom[10654] = 16'hfd8a;
  rom[10655] = 16'hfd89;
  rom[10656] = 16'hfd88;
  rom[10657] = 16'hfd86;
  rom[10658] = 16'hfd87;
  rom[10659] = 16'hfda8;
  rom[10660] = 16'hf588;
  rom[10661] = 16'hf5ca;
  rom[10662] = 16'hf5cc;
  rom[10663] = 16'hdd4c;
  rom[10664] = 16'hbc8b;
  rom[10665] = 16'h8307;
  rom[10666] = 16'h9c0e;
  rom[10667] = 16'he699;
  rom[10668] = 16'hffdf;
  rom[10669] = 16'hffff;
  rom[10670] = 16'hffff;
  rom[10671] = 16'hffff;
  rom[10672] = 16'hffff;
  rom[10673] = 16'hffff;
  rom[10674] = 16'hffff;
  rom[10675] = 16'hffff;
  rom[10676] = 16'hffff;
  rom[10677] = 16'hffff;
  rom[10678] = 16'hffff;
  rom[10679] = 16'hffff;
  rom[10680] = 16'hffff;
  rom[10681] = 16'hffff;
  rom[10682] = 16'hffff;
  rom[10683] = 16'hffff;
  rom[10684] = 16'hffff;
  rom[10685] = 16'hffff;
  rom[10686] = 16'hffff;
  rom[10687] = 16'hffff;
  rom[10688] = 16'hffde;
  rom[10689] = 16'hde98;
  rom[10690] = 16'haccf;
  rom[10691] = 16'h6aa6;
  rom[10692] = 16'hb4cd;
  rom[10693] = 16'hddee;
  rom[10694] = 16'hee2c;
  rom[10695] = 16'hf669;
  rom[10696] = 16'hf648;
  rom[10697] = 16'hee48;
  rom[10698] = 16'hee6a;
  rom[10699] = 16'hee6c;
  rom[10700] = 16'he60c;
  rom[10701] = 16'hcd8c;
  rom[10702] = 16'h7b46;
  rom[10703] = 16'h7b27;
  rom[10704] = 16'hc592;
  rom[10705] = 16'hf75a;
  rom[10706] = 16'hffff;
  rom[10707] = 16'hffdf;
  rom[10708] = 16'hffff;
  rom[10709] = 16'hffff;
  rom[10710] = 16'hffff;
  rom[10711] = 16'hffff;
  rom[10712] = 16'hffff;
  rom[10713] = 16'hffff;
  rom[10714] = 16'hffff;
  rom[10715] = 16'hffff;
  rom[10716] = 16'hffff;
  rom[10717] = 16'hffff;
  rom[10718] = 16'hffff;
  rom[10719] = 16'hffff;
  rom[10720] = 16'hffff;
  rom[10721] = 16'hffff;
  rom[10722] = 16'hffff;
  rom[10723] = 16'hffff;
  rom[10724] = 16'hffff;
  rom[10725] = 16'hf7df;
  rom[10726] = 16'hef7e;
  rom[10727] = 16'hb534;
  rom[10728] = 16'h7aea;
  rom[10729] = 16'h8b68;
  rom[10730] = 16'hd52d;
  rom[10731] = 16'hedcc;
  rom[10732] = 16'hfdca;
  rom[10733] = 16'hfda9;
  rom[10734] = 16'hf5a8;
  rom[10735] = 16'hf588;
  rom[10736] = 16'hfdc9;
  rom[10737] = 16'hfda8;
  rom[10738] = 16'hfd68;
  rom[10739] = 16'hfd69;
  rom[10740] = 16'hfd89;
  rom[10741] = 16'hfd48;
  rom[10742] = 16'hfd88;
  rom[10743] = 16'hfd68;
  rom[10744] = 16'hfd89;
  rom[10745] = 16'hf547;
  rom[10746] = 16'hfd89;
  rom[10747] = 16'hed2a;
  rom[10748] = 16'hd50c;
  rom[10749] = 16'h7b48;
  rom[10750] = 16'hffbe;
  rom[10751] = 16'hce59;
  rom[10752] = 16'h6aea;
  rom[10753] = 16'h6aa9;
  rom[10754] = 16'heefa;
  rom[10755] = 16'hffff;
  rom[10756] = 16'hffff;
  rom[10757] = 16'hffdf;
  rom[10758] = 16'hffff;
  rom[10759] = 16'hffff;
  rom[10760] = 16'hffff;
  rom[10761] = 16'hffff;
  rom[10762] = 16'hffff;
  rom[10763] = 16'hffff;
  rom[10764] = 16'hffff;
  rom[10765] = 16'hffff;
  rom[10766] = 16'hffff;
  rom[10767] = 16'hffff;
  rom[10768] = 16'hffff;
  rom[10769] = 16'hffff;
  rom[10770] = 16'hffff;
  rom[10771] = 16'hffff;
  rom[10772] = 16'hffff;
  rom[10773] = 16'hffff;
  rom[10774] = 16'hffff;
  rom[10775] = 16'hffff;
  rom[10776] = 16'hffff;
  rom[10777] = 16'hffff;
  rom[10778] = 16'hffff;
  rom[10779] = 16'hffff;
  rom[10780] = 16'hffff;
  rom[10781] = 16'hffff;
  rom[10782] = 16'hffff;
  rom[10783] = 16'hffff;
  rom[10784] = 16'hffff;
  rom[10785] = 16'hffff;
  rom[10786] = 16'hffff;
  rom[10787] = 16'hffff;
  rom[10788] = 16'hffff;
  rom[10789] = 16'hffff;
  rom[10790] = 16'hffff;
  rom[10791] = 16'hffff;
  rom[10792] = 16'hffff;
  rom[10793] = 16'hffff;
  rom[10794] = 16'hffff;
  rom[10795] = 16'hffff;
  rom[10796] = 16'hffff;
  rom[10797] = 16'hffff;
  rom[10798] = 16'hffff;
  rom[10799] = 16'hffff;
  rom[10800] = 16'hffff;
  rom[10801] = 16'hffff;
  rom[10802] = 16'hffff;
  rom[10803] = 16'hffff;
  rom[10804] = 16'hffff;
  rom[10805] = 16'hffff;
  rom[10806] = 16'hffff;
  rom[10807] = 16'hffff;
  rom[10808] = 16'hffff;
  rom[10809] = 16'hffff;
  rom[10810] = 16'hffff;
  rom[10811] = 16'hffff;
  rom[10812] = 16'hffff;
  rom[10813] = 16'hffff;
  rom[10814] = 16'hffff;
  rom[10815] = 16'hffff;
  rom[10816] = 16'hffff;
  rom[10817] = 16'hffff;
  rom[10818] = 16'hffff;
  rom[10819] = 16'hffff;
  rom[10820] = 16'hffff;
  rom[10821] = 16'hffff;
  rom[10822] = 16'hffff;
  rom[10823] = 16'hffff;
  rom[10824] = 16'hffff;
  rom[10825] = 16'hffff;
  rom[10826] = 16'hffff;
  rom[10827] = 16'hffff;
  rom[10828] = 16'hffff;
  rom[10829] = 16'hffff;
  rom[10830] = 16'hffff;
  rom[10831] = 16'hffff;
  rom[10832] = 16'hffff;
  rom[10833] = 16'hffff;
  rom[10834] = 16'hffff;
  rom[10835] = 16'hffff;
  rom[10836] = 16'hffdf;
  rom[10837] = 16'hffff;
  rom[10838] = 16'hffff;
  rom[10839] = 16'hffff;
  rom[10840] = 16'hffdf;
  rom[10841] = 16'hffff;
  rom[10842] = 16'hffde;
  rom[10843] = 16'hfffe;
  rom[10844] = 16'hb4ef;
  rom[10845] = 16'ha3c8;
  rom[10846] = 16'he52b;
  rom[10847] = 16'hfd6a;
  rom[10848] = 16'hfd48;
  rom[10849] = 16'hfd48;
  rom[10850] = 16'hf548;
  rom[10851] = 16'hfd68;
  rom[10852] = 16'hfd68;
  rom[10853] = 16'hfd69;
  rom[10854] = 16'hf568;
  rom[10855] = 16'hfda9;
  rom[10856] = 16'hfd67;
  rom[10857] = 16'hfda7;
  rom[10858] = 16'hf587;
  rom[10859] = 16'hfdc9;
  rom[10860] = 16'he569;
  rom[10861] = 16'hedcd;
  rom[10862] = 16'hdd8e;
  rom[10863] = 16'h82e5;
  rom[10864] = 16'h93ab;
  rom[10865] = 16'hde16;
  rom[10866] = 16'hff9c;
  rom[10867] = 16'hffff;
  rom[10868] = 16'hffff;
  rom[10869] = 16'hffff;
  rom[10870] = 16'hffff;
  rom[10871] = 16'hffff;
  rom[10872] = 16'hffff;
  rom[10873] = 16'hffff;
  rom[10874] = 16'hffff;
  rom[10875] = 16'hffff;
  rom[10876] = 16'hffff;
  rom[10877] = 16'hffff;
  rom[10878] = 16'hffff;
  rom[10879] = 16'hffff;
  rom[10880] = 16'hffff;
  rom[10881] = 16'hffff;
  rom[10882] = 16'hffff;
  rom[10883] = 16'hffff;
  rom[10884] = 16'hffff;
  rom[10885] = 16'hffff;
  rom[10886] = 16'hffbf;
  rom[10887] = 16'hffff;
  rom[10888] = 16'hffdf;
  rom[10889] = 16'hffff;
  rom[10890] = 16'hf77b;
  rom[10891] = 16'hde98;
  rom[10892] = 16'h8bec;
  rom[10893] = 16'h72e6;
  rom[10894] = 16'hc54c;
  rom[10895] = 16'he64d;
  rom[10896] = 16'hee4b;
  rom[10897] = 16'hee6b;
  rom[10898] = 16'heead;
  rom[10899] = 16'hd5ec;
  rom[10900] = 16'h9c28;
  rom[10901] = 16'h6b06;
  rom[10902] = 16'hb571;
  rom[10903] = 16'hf75a;
  rom[10904] = 16'hffbd;
  rom[10905] = 16'hffff;
  rom[10906] = 16'hffdf;
  rom[10907] = 16'hffff;
  rom[10908] = 16'hffdf;
  rom[10909] = 16'hffff;
  rom[10910] = 16'hffff;
  rom[10911] = 16'hffff;
  rom[10912] = 16'hffff;
  rom[10913] = 16'hffff;
  rom[10914] = 16'hffff;
  rom[10915] = 16'hffff;
  rom[10916] = 16'hffff;
  rom[10917] = 16'hffff;
  rom[10918] = 16'hffff;
  rom[10919] = 16'hffff;
  rom[10920] = 16'hffff;
  rom[10921] = 16'hffff;
  rom[10922] = 16'hffff;
  rom[10923] = 16'hffff;
  rom[10924] = 16'hffff;
  rom[10925] = 16'hffff;
  rom[10926] = 16'hffff;
  rom[10927] = 16'hffbf;
  rom[10928] = 16'heefb;
  rom[10929] = 16'hbcf1;
  rom[10930] = 16'h72e7;
  rom[10931] = 16'h93a7;
  rom[10932] = 16'he58d;
  rom[10933] = 16'hf5ab;
  rom[10934] = 16'hed69;
  rom[10935] = 16'hfda9;
  rom[10936] = 16'hfd68;
  rom[10937] = 16'hfd88;
  rom[10938] = 16'hfd68;
  rom[10939] = 16'hfd69;
  rom[10940] = 16'hfd69;
  rom[10941] = 16'hfd67;
  rom[10942] = 16'hf547;
  rom[10943] = 16'hfd88;
  rom[10944] = 16'hfd48;
  rom[10945] = 16'hfd67;
  rom[10946] = 16'hf547;
  rom[10947] = 16'hfd69;
  rom[10948] = 16'hdd2b;
  rom[10949] = 16'h8b68;
  rom[10950] = 16'hc5d4;
  rom[10951] = 16'hce16;
  rom[10952] = 16'h7b2a;
  rom[10953] = 16'h7ae9;
  rom[10954] = 16'hd636;
  rom[10955] = 16'hffff;
  rom[10956] = 16'hffff;
  rom[10957] = 16'hffff;
  rom[10958] = 16'hffdf;
  rom[10959] = 16'hffff;
  rom[10960] = 16'hffff;
  rom[10961] = 16'hffff;
  rom[10962] = 16'hffff;
  rom[10963] = 16'hffff;
  rom[10964] = 16'hffff;
  rom[10965] = 16'hffff;
  rom[10966] = 16'hffff;
  rom[10967] = 16'hffff;
  rom[10968] = 16'hffff;
  rom[10969] = 16'hffff;
  rom[10970] = 16'hffff;
  rom[10971] = 16'hffff;
  rom[10972] = 16'hffff;
  rom[10973] = 16'hffff;
  rom[10974] = 16'hffff;
  rom[10975] = 16'hffff;
  rom[10976] = 16'hffff;
  rom[10977] = 16'hffff;
  rom[10978] = 16'hffff;
  rom[10979] = 16'hffff;
  rom[10980] = 16'hffff;
  rom[10981] = 16'hffff;
  rom[10982] = 16'hffff;
  rom[10983] = 16'hffff;
  rom[10984] = 16'hffff;
  rom[10985] = 16'hffff;
  rom[10986] = 16'hffff;
  rom[10987] = 16'hffff;
  rom[10988] = 16'hffff;
  rom[10989] = 16'hffff;
  rom[10990] = 16'hffff;
  rom[10991] = 16'hffff;
  rom[10992] = 16'hffff;
  rom[10993] = 16'hffff;
  rom[10994] = 16'hffff;
  rom[10995] = 16'hffff;
  rom[10996] = 16'hffff;
  rom[10997] = 16'hffff;
  rom[10998] = 16'hffff;
  rom[10999] = 16'hffff;
  rom[11000] = 16'hffff;
  rom[11001] = 16'hffff;
  rom[11002] = 16'hffff;
  rom[11003] = 16'hffff;
  rom[11004] = 16'hffff;
  rom[11005] = 16'hffff;
  rom[11006] = 16'hffff;
  rom[11007] = 16'hffff;
  rom[11008] = 16'hffff;
  rom[11009] = 16'hffff;
  rom[11010] = 16'hffff;
  rom[11011] = 16'hffff;
  rom[11012] = 16'hffff;
  rom[11013] = 16'hffff;
  rom[11014] = 16'hffff;
  rom[11015] = 16'hffff;
  rom[11016] = 16'hffff;
  rom[11017] = 16'hffff;
  rom[11018] = 16'hffff;
  rom[11019] = 16'hffff;
  rom[11020] = 16'hffff;
  rom[11021] = 16'hffff;
  rom[11022] = 16'hffff;
  rom[11023] = 16'hffff;
  rom[11024] = 16'hffff;
  rom[11025] = 16'hffff;
  rom[11026] = 16'hffff;
  rom[11027] = 16'hffff;
  rom[11028] = 16'hffff;
  rom[11029] = 16'hffff;
  rom[11030] = 16'hffff;
  rom[11031] = 16'hffff;
  rom[11032] = 16'hffff;
  rom[11033] = 16'hffff;
  rom[11034] = 16'hffff;
  rom[11035] = 16'hffff;
  rom[11036] = 16'hffff;
  rom[11037] = 16'hffff;
  rom[11038] = 16'hffff;
  rom[11039] = 16'hffdf;
  rom[11040] = 16'hffff;
  rom[11041] = 16'hffdf;
  rom[11042] = 16'hffff;
  rom[11043] = 16'hff9c;
  rom[11044] = 16'h9c0c;
  rom[11045] = 16'hcd0c;
  rom[11046] = 16'hed6b;
  rom[11047] = 16'hf528;
  rom[11048] = 16'hfd48;
  rom[11049] = 16'hfd48;
  rom[11050] = 16'hfd69;
  rom[11051] = 16'hfd68;
  rom[11052] = 16'hfd89;
  rom[11053] = 16'hfd67;
  rom[11054] = 16'hfd88;
  rom[11055] = 16'hfd89;
  rom[11056] = 16'hfd89;
  rom[11057] = 16'hfda8;
  rom[11058] = 16'hf589;
  rom[11059] = 16'hedab;
  rom[11060] = 16'he5ed;
  rom[11061] = 16'hbd0c;
  rom[11062] = 16'h5a03;
  rom[11063] = 16'hb4f0;
  rom[11064] = 16'hff5b;
  rom[11065] = 16'hffde;
  rom[11066] = 16'hffff;
  rom[11067] = 16'hffff;
  rom[11068] = 16'hffff;
  rom[11069] = 16'hffff;
  rom[11070] = 16'hffff;
  rom[11071] = 16'hffff;
  rom[11072] = 16'hffff;
  rom[11073] = 16'hffff;
  rom[11074] = 16'hffff;
  rom[11075] = 16'hffff;
  rom[11076] = 16'hffff;
  rom[11077] = 16'hffdf;
  rom[11078] = 16'hffff;
  rom[11079] = 16'hffff;
  rom[11080] = 16'hffff;
  rom[11081] = 16'hffff;
  rom[11082] = 16'hffff;
  rom[11083] = 16'hffff;
  rom[11084] = 16'hffff;
  rom[11085] = 16'hffff;
  rom[11086] = 16'hffff;
  rom[11087] = 16'hffff;
  rom[11088] = 16'hffbf;
  rom[11089] = 16'hffff;
  rom[11090] = 16'hffff;
  rom[11091] = 16'hfffe;
  rom[11092] = 16'hff9d;
  rom[11093] = 16'hbd53;
  rom[11094] = 16'h6285;
  rom[11095] = 16'hc54d;
  rom[11096] = 16'he64f;
  rom[11097] = 16'he64f;
  rom[11098] = 16'hd60e;
  rom[11099] = 16'h8387;
  rom[11100] = 16'h7b28;
  rom[11101] = 16'he6d9;
  rom[11102] = 16'hffff;
  rom[11103] = 16'hffff;
  rom[11104] = 16'hffff;
  rom[11105] = 16'hffff;
  rom[11106] = 16'hffff;
  rom[11107] = 16'hffff;
  rom[11108] = 16'hffff;
  rom[11109] = 16'hffdf;
  rom[11110] = 16'hffff;
  rom[11111] = 16'hffdf;
  rom[11112] = 16'hffff;
  rom[11113] = 16'hffff;
  rom[11114] = 16'hffff;
  rom[11115] = 16'hffff;
  rom[11116] = 16'hffff;
  rom[11117] = 16'hffff;
  rom[11118] = 16'hffff;
  rom[11119] = 16'hffff;
  rom[11120] = 16'hffff;
  rom[11121] = 16'hffff;
  rom[11122] = 16'hffff;
  rom[11123] = 16'hffff;
  rom[11124] = 16'hffff;
  rom[11125] = 16'hffde;
  rom[11126] = 16'hffff;
  rom[11127] = 16'hffff;
  rom[11128] = 16'hffff;
  rom[11129] = 16'hffdf;
  rom[11130] = 16'he6b9;
  rom[11131] = 16'h72e8;
  rom[11132] = 16'h8b47;
  rom[11133] = 16'hdd6c;
  rom[11134] = 16'hf5cd;
  rom[11135] = 16'hf569;
  rom[11136] = 16'hf568;
  rom[11137] = 16'hfd88;
  rom[11138] = 16'hfd89;
  rom[11139] = 16'hfd69;
  rom[11140] = 16'hfd69;
  rom[11141] = 16'hfd88;
  rom[11142] = 16'hfd67;
  rom[11143] = 16'hfd68;
  rom[11144] = 16'hfd69;
  rom[11145] = 16'hfd68;
  rom[11146] = 16'hfd67;
  rom[11147] = 16'hf527;
  rom[11148] = 16'hed0a;
  rom[11149] = 16'hac29;
  rom[11150] = 16'h9c4e;
  rom[11151] = 16'hc5d5;
  rom[11152] = 16'h832a;
  rom[11153] = 16'h93ab;
  rom[11154] = 16'hcdd5;
  rom[11155] = 16'hffff;
  rom[11156] = 16'hffff;
  rom[11157] = 16'hffff;
  rom[11158] = 16'hffff;
  rom[11159] = 16'hffff;
  rom[11160] = 16'hffff;
  rom[11161] = 16'hffff;
  rom[11162] = 16'hffff;
  rom[11163] = 16'hffff;
  rom[11164] = 16'hffff;
  rom[11165] = 16'hffff;
  rom[11166] = 16'hffff;
  rom[11167] = 16'hffff;
  rom[11168] = 16'hffff;
  rom[11169] = 16'hffff;
  rom[11170] = 16'hffff;
  rom[11171] = 16'hffff;
  rom[11172] = 16'hffff;
  rom[11173] = 16'hffff;
  rom[11174] = 16'hffff;
  rom[11175] = 16'hffff;
  rom[11176] = 16'hffff;
  rom[11177] = 16'hffff;
  rom[11178] = 16'hffff;
  rom[11179] = 16'hffff;
  rom[11180] = 16'hffff;
  rom[11181] = 16'hffff;
  rom[11182] = 16'hffff;
  rom[11183] = 16'hffff;
  rom[11184] = 16'hffff;
  rom[11185] = 16'hffff;
  rom[11186] = 16'hffff;
  rom[11187] = 16'hffff;
  rom[11188] = 16'hffff;
  rom[11189] = 16'hffff;
  rom[11190] = 16'hffff;
  rom[11191] = 16'hffff;
  rom[11192] = 16'hffff;
  rom[11193] = 16'hffff;
  rom[11194] = 16'hffff;
  rom[11195] = 16'hffff;
  rom[11196] = 16'hffff;
  rom[11197] = 16'hffff;
  rom[11198] = 16'hffff;
  rom[11199] = 16'hffff;
  rom[11200] = 16'hffff;
  rom[11201] = 16'hffff;
  rom[11202] = 16'hffff;
  rom[11203] = 16'hffff;
  rom[11204] = 16'hffff;
  rom[11205] = 16'hffff;
  rom[11206] = 16'hffff;
  rom[11207] = 16'hffff;
  rom[11208] = 16'hffff;
  rom[11209] = 16'hffff;
  rom[11210] = 16'hffff;
  rom[11211] = 16'hffff;
  rom[11212] = 16'hffff;
  rom[11213] = 16'hffff;
  rom[11214] = 16'hffff;
  rom[11215] = 16'hffff;
  rom[11216] = 16'hffff;
  rom[11217] = 16'hffff;
  rom[11218] = 16'hffff;
  rom[11219] = 16'hffff;
  rom[11220] = 16'hffff;
  rom[11221] = 16'hffff;
  rom[11222] = 16'hffff;
  rom[11223] = 16'hffff;
  rom[11224] = 16'hffff;
  rom[11225] = 16'hffff;
  rom[11226] = 16'hffff;
  rom[11227] = 16'hffff;
  rom[11228] = 16'hffff;
  rom[11229] = 16'hffff;
  rom[11230] = 16'hffff;
  rom[11231] = 16'hffff;
  rom[11232] = 16'hffff;
  rom[11233] = 16'hffff;
  rom[11234] = 16'hffff;
  rom[11235] = 16'hffff;
  rom[11236] = 16'hffff;
  rom[11237] = 16'hffff;
  rom[11238] = 16'hffff;
  rom[11239] = 16'hffff;
  rom[11240] = 16'hffff;
  rom[11241] = 16'hffff;
  rom[11242] = 16'hffff;
  rom[11243] = 16'heeb8;
  rom[11244] = 16'h8b47;
  rom[11245] = 16'hdd4b;
  rom[11246] = 16'hed28;
  rom[11247] = 16'hfd49;
  rom[11248] = 16'hfd47;
  rom[11249] = 16'hfd48;
  rom[11250] = 16'hfd68;
  rom[11251] = 16'hf589;
  rom[11252] = 16'hf588;
  rom[11253] = 16'hfd47;
  rom[11254] = 16'hfd67;
  rom[11255] = 16'hfd88;
  rom[11256] = 16'hfd68;
  rom[11257] = 16'hfd89;
  rom[11258] = 16'hedab;
  rom[11259] = 16'he5cd;
  rom[11260] = 16'h9c29;
  rom[11261] = 16'h7b48;
  rom[11262] = 16'hd635;
  rom[11263] = 16'hffbd;
  rom[11264] = 16'hfffe;
  rom[11265] = 16'hffff;
  rom[11266] = 16'hffff;
  rom[11267] = 16'hffff;
  rom[11268] = 16'hffff;
  rom[11269] = 16'hffff;
  rom[11270] = 16'hffff;
  rom[11271] = 16'hffff;
  rom[11272] = 16'hffff;
  rom[11273] = 16'hffff;
  rom[11274] = 16'hffff;
  rom[11275] = 16'hffff;
  rom[11276] = 16'hffff;
  rom[11277] = 16'hffff;
  rom[11278] = 16'hffff;
  rom[11279] = 16'hffff;
  rom[11280] = 16'hffff;
  rom[11281] = 16'hffff;
  rom[11282] = 16'hffff;
  rom[11283] = 16'hffff;
  rom[11284] = 16'hffff;
  rom[11285] = 16'hffff;
  rom[11286] = 16'hffff;
  rom[11287] = 16'hffff;
  rom[11288] = 16'hffff;
  rom[11289] = 16'hffff;
  rom[11290] = 16'hffff;
  rom[11291] = 16'hffff;
  rom[11292] = 16'hffff;
  rom[11293] = 16'hffde;
  rom[11294] = 16'hd636;
  rom[11295] = 16'h7b49;
  rom[11296] = 16'h942b;
  rom[11297] = 16'hbd4f;
  rom[11298] = 16'h7347;
  rom[11299] = 16'ha4cf;
  rom[11300] = 16'hf77b;
  rom[11301] = 16'hffff;
  rom[11302] = 16'hffdf;
  rom[11303] = 16'hffff;
  rom[11304] = 16'hffff;
  rom[11305] = 16'hffff;
  rom[11306] = 16'hffff;
  rom[11307] = 16'hffff;
  rom[11308] = 16'hffff;
  rom[11309] = 16'hffff;
  rom[11310] = 16'hffff;
  rom[11311] = 16'hffff;
  rom[11312] = 16'hffff;
  rom[11313] = 16'hffff;
  rom[11314] = 16'hffff;
  rom[11315] = 16'hffff;
  rom[11316] = 16'hffff;
  rom[11317] = 16'hffff;
  rom[11318] = 16'hffff;
  rom[11319] = 16'hffff;
  rom[11320] = 16'hffff;
  rom[11321] = 16'hffff;
  rom[11322] = 16'hffff;
  rom[11323] = 16'hffff;
  rom[11324] = 16'hffff;
  rom[11325] = 16'hffff;
  rom[11326] = 16'hffde;
  rom[11327] = 16'hffff;
  rom[11328] = 16'hffff;
  rom[11329] = 16'hffff;
  rom[11330] = 16'hffff;
  rom[11331] = 16'hff7d;
  rom[11332] = 16'h942e;
  rom[11333] = 16'h8327;
  rom[11334] = 16'hcd2d;
  rom[11335] = 16'hed6c;
  rom[11336] = 16'hf5ca;
  rom[11337] = 16'hfd89;
  rom[11338] = 16'hfd67;
  rom[11339] = 16'hfd68;
  rom[11340] = 16'hfd67;
  rom[11341] = 16'hfd68;
  rom[11342] = 16'hf568;
  rom[11343] = 16'hfd6a;
  rom[11344] = 16'hf549;
  rom[11345] = 16'hfd68;
  rom[11346] = 16'hfd47;
  rom[11347] = 16'hfd68;
  rom[11348] = 16'hf569;
  rom[11349] = 16'hc4aa;
  rom[11350] = 16'h6285;
  rom[11351] = 16'ha46e;
  rom[11352] = 16'h8348;
  rom[11353] = 16'hac4d;
  rom[11354] = 16'hb4d1;
  rom[11355] = 16'hffff;
  rom[11356] = 16'hf7ff;
  rom[11357] = 16'hffff;
  rom[11358] = 16'hffdf;
  rom[11359] = 16'hffff;
  rom[11360] = 16'hffff;
  rom[11361] = 16'hffff;
  rom[11362] = 16'hffff;
  rom[11363] = 16'hffff;
  rom[11364] = 16'hffff;
  rom[11365] = 16'hffff;
  rom[11366] = 16'hffff;
  rom[11367] = 16'hffff;
  rom[11368] = 16'hffff;
  rom[11369] = 16'hffff;
  rom[11370] = 16'hffff;
  rom[11371] = 16'hffff;
  rom[11372] = 16'hffff;
  rom[11373] = 16'hffff;
  rom[11374] = 16'hffff;
  rom[11375] = 16'hffff;
  rom[11376] = 16'hffff;
  rom[11377] = 16'hffff;
  rom[11378] = 16'hffff;
  rom[11379] = 16'hffff;
  rom[11380] = 16'hffff;
  rom[11381] = 16'hffff;
  rom[11382] = 16'hffff;
  rom[11383] = 16'hffff;
  rom[11384] = 16'hffff;
  rom[11385] = 16'hffff;
  rom[11386] = 16'hffff;
  rom[11387] = 16'hffff;
  rom[11388] = 16'hffff;
  rom[11389] = 16'hffff;
  rom[11390] = 16'hffff;
  rom[11391] = 16'hffff;
  rom[11392] = 16'hffff;
  rom[11393] = 16'hffff;
  rom[11394] = 16'hffff;
  rom[11395] = 16'hffff;
  rom[11396] = 16'hffff;
  rom[11397] = 16'hffff;
  rom[11398] = 16'hffff;
  rom[11399] = 16'hffff;
  rom[11400] = 16'hffff;
  rom[11401] = 16'hffff;
  rom[11402] = 16'hffff;
  rom[11403] = 16'hffff;
  rom[11404] = 16'hffff;
  rom[11405] = 16'hffff;
  rom[11406] = 16'hffff;
  rom[11407] = 16'hffff;
  rom[11408] = 16'hffff;
  rom[11409] = 16'hffff;
  rom[11410] = 16'hffff;
  rom[11411] = 16'hffff;
  rom[11412] = 16'hffff;
  rom[11413] = 16'hffff;
  rom[11414] = 16'hffff;
  rom[11415] = 16'hffff;
  rom[11416] = 16'hffff;
  rom[11417] = 16'hffff;
  rom[11418] = 16'hffff;
  rom[11419] = 16'hffff;
  rom[11420] = 16'hffff;
  rom[11421] = 16'hffff;
  rom[11422] = 16'hffff;
  rom[11423] = 16'hffff;
  rom[11424] = 16'hffff;
  rom[11425] = 16'hffff;
  rom[11426] = 16'hffff;
  rom[11427] = 16'hffff;
  rom[11428] = 16'hffff;
  rom[11429] = 16'hffff;
  rom[11430] = 16'hffff;
  rom[11431] = 16'hffff;
  rom[11432] = 16'hffff;
  rom[11433] = 16'hffff;
  rom[11434] = 16'hffff;
  rom[11435] = 16'hffbf;
  rom[11436] = 16'hffff;
  rom[11437] = 16'hffff;
  rom[11438] = 16'hef7d;
  rom[11439] = 16'hffff;
  rom[11440] = 16'hffdf;
  rom[11441] = 16'hffff;
  rom[11442] = 16'hffff;
  rom[11443] = 16'hcdd4;
  rom[11444] = 16'ha3c9;
  rom[11445] = 16'he54b;
  rom[11446] = 16'hfd89;
  rom[11447] = 16'hfd68;
  rom[11448] = 16'hfd49;
  rom[11449] = 16'hfd49;
  rom[11450] = 16'hf56a;
  rom[11451] = 16'hed69;
  rom[11452] = 16'hfda9;
  rom[11453] = 16'hfd87;
  rom[11454] = 16'hfd67;
  rom[11455] = 16'hfd68;
  rom[11456] = 16'hfd89;
  rom[11457] = 16'hf56a;
  rom[11458] = 16'hed8d;
  rom[11459] = 16'h8b87;
  rom[11460] = 16'h6ae7;
  rom[11461] = 16'hdeb8;
  rom[11462] = 16'hfffe;
  rom[11463] = 16'hffff;
  rom[11464] = 16'hffff;
  rom[11465] = 16'hffff;
  rom[11466] = 16'hffff;
  rom[11467] = 16'hffff;
  rom[11468] = 16'hffff;
  rom[11469] = 16'hffff;
  rom[11470] = 16'hffff;
  rom[11471] = 16'hffff;
  rom[11472] = 16'hffff;
  rom[11473] = 16'hffff;
  rom[11474] = 16'hffff;
  rom[11475] = 16'hffff;
  rom[11476] = 16'hffff;
  rom[11477] = 16'hffff;
  rom[11478] = 16'hffff;
  rom[11479] = 16'hffff;
  rom[11480] = 16'hffff;
  rom[11481] = 16'hffff;
  rom[11482] = 16'hffff;
  rom[11483] = 16'hffff;
  rom[11484] = 16'hffff;
  rom[11485] = 16'hffff;
  rom[11486] = 16'hffff;
  rom[11487] = 16'hffff;
  rom[11488] = 16'hffff;
  rom[11489] = 16'hffff;
  rom[11490] = 16'hffff;
  rom[11491] = 16'hffff;
  rom[11492] = 16'hffff;
  rom[11493] = 16'hffff;
  rom[11494] = 16'hffff;
  rom[11495] = 16'he6f9;
  rom[11496] = 16'h83ac;
  rom[11497] = 16'h3983;
  rom[11498] = 16'hbd73;
  rom[11499] = 16'hff9c;
  rom[11500] = 16'hffff;
  rom[11501] = 16'hffdf;
  rom[11502] = 16'hffff;
  rom[11503] = 16'hffff;
  rom[11504] = 16'hffff;
  rom[11505] = 16'hffff;
  rom[11506] = 16'hffff;
  rom[11507] = 16'hffff;
  rom[11508] = 16'hffff;
  rom[11509] = 16'hffff;
  rom[11510] = 16'hffff;
  rom[11511] = 16'hffff;
  rom[11512] = 16'hffff;
  rom[11513] = 16'hffff;
  rom[11514] = 16'hffff;
  rom[11515] = 16'hffff;
  rom[11516] = 16'hffff;
  rom[11517] = 16'hffff;
  rom[11518] = 16'hffff;
  rom[11519] = 16'hffff;
  rom[11520] = 16'hffff;
  rom[11521] = 16'hffff;
  rom[11522] = 16'hffff;
  rom[11523] = 16'hffff;
  rom[11524] = 16'hffff;
  rom[11525] = 16'hffdf;
  rom[11526] = 16'hffbf;
  rom[11527] = 16'hffbd;
  rom[11528] = 16'hffff;
  rom[11529] = 16'hffff;
  rom[11530] = 16'hffff;
  rom[11531] = 16'hffff;
  rom[11532] = 16'hfffe;
  rom[11533] = 16'ha4af;
  rom[11534] = 16'h72c5;
  rom[11535] = 16'hd52d;
  rom[11536] = 16'hed8c;
  rom[11537] = 16'hed49;
  rom[11538] = 16'hfd88;
  rom[11539] = 16'hfd67;
  rom[11540] = 16'hfd87;
  rom[11541] = 16'hfd68;
  rom[11542] = 16'hfd8a;
  rom[11543] = 16'hf56a;
  rom[11544] = 16'hfd6a;
  rom[11545] = 16'hfd48;
  rom[11546] = 16'hfd48;
  rom[11547] = 16'hfd48;
  rom[11548] = 16'hed08;
  rom[11549] = 16'hd52c;
  rom[11550] = 16'h9389;
  rom[11551] = 16'h8348;
  rom[11552] = 16'ha40a;
  rom[11553] = 16'hac2c;
  rom[11554] = 16'ha3ee;
  rom[11555] = 16'hffdf;
  rom[11556] = 16'hffff;
  rom[11557] = 16'hf7ff;
  rom[11558] = 16'hffff;
  rom[11559] = 16'hffff;
  rom[11560] = 16'hffff;
  rom[11561] = 16'hffff;
  rom[11562] = 16'hffff;
  rom[11563] = 16'hffff;
  rom[11564] = 16'hffff;
  rom[11565] = 16'hffff;
  rom[11566] = 16'hffff;
  rom[11567] = 16'hffff;
  rom[11568] = 16'hffff;
  rom[11569] = 16'hffff;
  rom[11570] = 16'hffff;
  rom[11571] = 16'hffff;
  rom[11572] = 16'hffff;
  rom[11573] = 16'hffff;
  rom[11574] = 16'hffff;
  rom[11575] = 16'hffff;
  rom[11576] = 16'hffff;
  rom[11577] = 16'hffff;
  rom[11578] = 16'hffff;
  rom[11579] = 16'hffff;
  rom[11580] = 16'hffff;
  rom[11581] = 16'hffff;
  rom[11582] = 16'hffff;
  rom[11583] = 16'hffff;
  rom[11584] = 16'hffff;
  rom[11585] = 16'hffff;
  rom[11586] = 16'hffff;
  rom[11587] = 16'hffff;
  rom[11588] = 16'hffff;
  rom[11589] = 16'hffff;
  rom[11590] = 16'hffff;
  rom[11591] = 16'hffff;
  rom[11592] = 16'hffff;
  rom[11593] = 16'hffff;
  rom[11594] = 16'hffff;
  rom[11595] = 16'hffff;
  rom[11596] = 16'hffff;
  rom[11597] = 16'hffff;
  rom[11598] = 16'hffff;
  rom[11599] = 16'hffff;
  rom[11600] = 16'hffff;
  rom[11601] = 16'hffff;
  rom[11602] = 16'hffff;
  rom[11603] = 16'hffff;
  rom[11604] = 16'hffff;
  rom[11605] = 16'hffff;
  rom[11606] = 16'hffff;
  rom[11607] = 16'hffff;
  rom[11608] = 16'hffff;
  rom[11609] = 16'hffff;
  rom[11610] = 16'hffff;
  rom[11611] = 16'hffff;
  rom[11612] = 16'hffff;
  rom[11613] = 16'hffff;
  rom[11614] = 16'hffff;
  rom[11615] = 16'hffff;
  rom[11616] = 16'hffff;
  rom[11617] = 16'hffff;
  rom[11618] = 16'hffff;
  rom[11619] = 16'hffff;
  rom[11620] = 16'hffff;
  rom[11621] = 16'hffff;
  rom[11622] = 16'hffff;
  rom[11623] = 16'hffff;
  rom[11624] = 16'hffff;
  rom[11625] = 16'hffff;
  rom[11626] = 16'hffff;
  rom[11627] = 16'hffff;
  rom[11628] = 16'hffff;
  rom[11629] = 16'hffff;
  rom[11630] = 16'hffff;
  rom[11631] = 16'hffff;
  rom[11632] = 16'hffff;
  rom[11633] = 16'hffff;
  rom[11634] = 16'hffff;
  rom[11635] = 16'hffff;
  rom[11636] = 16'hffdf;
  rom[11637] = 16'hffff;
  rom[11638] = 16'h844f;
  rom[11639] = 16'had33;
  rom[11640] = 16'hf79d;
  rom[11641] = 16'hffdf;
  rom[11642] = 16'hfffe;
  rom[11643] = 16'hb511;
  rom[11644] = 16'ha3c8;
  rom[11645] = 16'he52a;
  rom[11646] = 16'hf548;
  rom[11647] = 16'hfd47;
  rom[11648] = 16'hfd27;
  rom[11649] = 16'hfd69;
  rom[11650] = 16'hed49;
  rom[11651] = 16'hf589;
  rom[11652] = 16'hf588;
  rom[11653] = 16'hfd67;
  rom[11654] = 16'hf567;
  rom[11655] = 16'hfdc9;
  rom[11656] = 16'hed6a;
  rom[11657] = 16'hf5ae;
  rom[11658] = 16'hac09;
  rom[11659] = 16'h8348;
  rom[11660] = 16'hde77;
  rom[11661] = 16'hffdf;
  rom[11662] = 16'hffff;
  rom[11663] = 16'hffff;
  rom[11664] = 16'hffff;
  rom[11665] = 16'hffff;
  rom[11666] = 16'hffff;
  rom[11667] = 16'hffff;
  rom[11668] = 16'hffff;
  rom[11669] = 16'hffff;
  rom[11670] = 16'hffff;
  rom[11671] = 16'hffff;
  rom[11672] = 16'hffff;
  rom[11673] = 16'hffff;
  rom[11674] = 16'hffff;
  rom[11675] = 16'hffff;
  rom[11676] = 16'hffff;
  rom[11677] = 16'hffff;
  rom[11678] = 16'hffff;
  rom[11679] = 16'hffff;
  rom[11680] = 16'hffff;
  rom[11681] = 16'hffff;
  rom[11682] = 16'hffff;
  rom[11683] = 16'hffff;
  rom[11684] = 16'hffff;
  rom[11685] = 16'hffff;
  rom[11686] = 16'hffff;
  rom[11687] = 16'hffff;
  rom[11688] = 16'hffff;
  rom[11689] = 16'hffff;
  rom[11690] = 16'hffff;
  rom[11691] = 16'hffff;
  rom[11692] = 16'hffff;
  rom[11693] = 16'hffff;
  rom[11694] = 16'hfffe;
  rom[11695] = 16'hffff;
  rom[11696] = 16'he6fa;
  rom[11697] = 16'he6b9;
  rom[11698] = 16'hffbd;
  rom[11699] = 16'hffff;
  rom[11700] = 16'hffff;
  rom[11701] = 16'hffff;
  rom[11702] = 16'hffff;
  rom[11703] = 16'hffff;
  rom[11704] = 16'hffff;
  rom[11705] = 16'hffff;
  rom[11706] = 16'hffff;
  rom[11707] = 16'hffff;
  rom[11708] = 16'hffff;
  rom[11709] = 16'hffff;
  rom[11710] = 16'hffff;
  rom[11711] = 16'hffff;
  rom[11712] = 16'hffff;
  rom[11713] = 16'hffff;
  rom[11714] = 16'hffff;
  rom[11715] = 16'hffff;
  rom[11716] = 16'hffff;
  rom[11717] = 16'hffff;
  rom[11718] = 16'hffff;
  rom[11719] = 16'hffff;
  rom[11720] = 16'hffff;
  rom[11721] = 16'hffff;
  rom[11722] = 16'hffff;
  rom[11723] = 16'hffff;
  rom[11724] = 16'hffff;
  rom[11725] = 16'hffff;
  rom[11726] = 16'hffff;
  rom[11727] = 16'hfffe;
  rom[11728] = 16'hffff;
  rom[11729] = 16'hffff;
  rom[11730] = 16'hffdf;
  rom[11731] = 16'hffdf;
  rom[11732] = 16'hffde;
  rom[11733] = 16'hfffe;
  rom[11734] = 16'hb510;
  rom[11735] = 16'h8b67;
  rom[11736] = 16'hd52c;
  rom[11737] = 16'hf5cd;
  rom[11738] = 16'hed48;
  rom[11739] = 16'hfda8;
  rom[11740] = 16'hf547;
  rom[11741] = 16'hfd88;
  rom[11742] = 16'hf568;
  rom[11743] = 16'hf569;
  rom[11744] = 16'hfd68;
  rom[11745] = 16'hfd68;
  rom[11746] = 16'hfd47;
  rom[11747] = 16'hfd48;
  rom[11748] = 16'hf569;
  rom[11749] = 16'he52c;
  rom[11750] = 16'h9346;
  rom[11751] = 16'h6202;
  rom[11752] = 16'hac2a;
  rom[11753] = 16'hbc8d;
  rom[11754] = 16'h93ac;
  rom[11755] = 16'hff7e;
  rom[11756] = 16'hffdf;
  rom[11757] = 16'hffff;
  rom[11758] = 16'hffff;
  rom[11759] = 16'hffff;
  rom[11760] = 16'hffff;
  rom[11761] = 16'hffff;
  rom[11762] = 16'hffff;
  rom[11763] = 16'hffff;
  rom[11764] = 16'hffff;
  rom[11765] = 16'hffff;
  rom[11766] = 16'hffff;
  rom[11767] = 16'hffff;
  rom[11768] = 16'hffff;
  rom[11769] = 16'hffff;
  rom[11770] = 16'hffff;
  rom[11771] = 16'hffff;
  rom[11772] = 16'hffff;
  rom[11773] = 16'hffff;
  rom[11774] = 16'hffff;
  rom[11775] = 16'hffff;
  rom[11776] = 16'hffff;
  rom[11777] = 16'hffff;
  rom[11778] = 16'hffff;
  rom[11779] = 16'hffff;
  rom[11780] = 16'hffff;
  rom[11781] = 16'hffff;
  rom[11782] = 16'hffff;
  rom[11783] = 16'hffff;
  rom[11784] = 16'hffff;
  rom[11785] = 16'hffff;
  rom[11786] = 16'hffff;
  rom[11787] = 16'hffff;
  rom[11788] = 16'hffff;
  rom[11789] = 16'hffff;
  rom[11790] = 16'hffff;
  rom[11791] = 16'hffff;
  rom[11792] = 16'hffff;
  rom[11793] = 16'hffff;
  rom[11794] = 16'hffff;
  rom[11795] = 16'hffff;
  rom[11796] = 16'hffff;
  rom[11797] = 16'hffff;
  rom[11798] = 16'hffff;
  rom[11799] = 16'hffff;
  rom[11800] = 16'hffff;
  rom[11801] = 16'hffff;
  rom[11802] = 16'hffff;
  rom[11803] = 16'hffff;
  rom[11804] = 16'hffff;
  rom[11805] = 16'hffff;
  rom[11806] = 16'hffff;
  rom[11807] = 16'hffff;
  rom[11808] = 16'hffff;
  rom[11809] = 16'hffff;
  rom[11810] = 16'hffff;
  rom[11811] = 16'hffff;
  rom[11812] = 16'hffff;
  rom[11813] = 16'hffff;
  rom[11814] = 16'hffff;
  rom[11815] = 16'hffff;
  rom[11816] = 16'hffff;
  rom[11817] = 16'hffff;
  rom[11818] = 16'hffff;
  rom[11819] = 16'hffff;
  rom[11820] = 16'hffff;
  rom[11821] = 16'hffff;
  rom[11822] = 16'hffff;
  rom[11823] = 16'hffff;
  rom[11824] = 16'hffff;
  rom[11825] = 16'hffff;
  rom[11826] = 16'hffff;
  rom[11827] = 16'hffff;
  rom[11828] = 16'hffff;
  rom[11829] = 16'hffff;
  rom[11830] = 16'hffff;
  rom[11831] = 16'hffff;
  rom[11832] = 16'hffff;
  rom[11833] = 16'hffff;
  rom[11834] = 16'hffff;
  rom[11835] = 16'hffff;
  rom[11836] = 16'hffdf;
  rom[11837] = 16'hffff;
  rom[11838] = 16'hb594;
  rom[11839] = 16'h31a3;
  rom[11840] = 16'h8bcd;
  rom[11841] = 16'hde58;
  rom[11842] = 16'hff9c;
  rom[11843] = 16'hac8e;
  rom[11844] = 16'habc7;
  rom[11845] = 16'hed6a;
  rom[11846] = 16'hfd48;
  rom[11847] = 16'hfd47;
  rom[11848] = 16'hfd69;
  rom[11849] = 16'hf568;
  rom[11850] = 16'hfd8a;
  rom[11851] = 16'hfd69;
  rom[11852] = 16'hfd68;
  rom[11853] = 16'hfda8;
  rom[11854] = 16'hfd88;
  rom[11855] = 16'hf5c9;
  rom[11856] = 16'he58c;
  rom[11857] = 16'hb44b;
  rom[11858] = 16'h8b49;
  rom[11859] = 16'hde36;
  rom[11860] = 16'hffff;
  rom[11861] = 16'hffff;
  rom[11862] = 16'hffff;
  rom[11863] = 16'hffff;
  rom[11864] = 16'hffff;
  rom[11865] = 16'hffff;
  rom[11866] = 16'hffff;
  rom[11867] = 16'hffff;
  rom[11868] = 16'hffff;
  rom[11869] = 16'hffff;
  rom[11870] = 16'hffff;
  rom[11871] = 16'hffff;
  rom[11872] = 16'hffff;
  rom[11873] = 16'hffff;
  rom[11874] = 16'hffff;
  rom[11875] = 16'hffff;
  rom[11876] = 16'hffff;
  rom[11877] = 16'hffff;
  rom[11878] = 16'hffff;
  rom[11879] = 16'hffff;
  rom[11880] = 16'hffff;
  rom[11881] = 16'hffff;
  rom[11882] = 16'hffff;
  rom[11883] = 16'hffff;
  rom[11884] = 16'hffff;
  rom[11885] = 16'hffff;
  rom[11886] = 16'hffff;
  rom[11887] = 16'hffff;
  rom[11888] = 16'hffff;
  rom[11889] = 16'hffff;
  rom[11890] = 16'hffff;
  rom[11891] = 16'hffff;
  rom[11892] = 16'hffff;
  rom[11893] = 16'hffff;
  rom[11894] = 16'hffff;
  rom[11895] = 16'hffff;
  rom[11896] = 16'hffff;
  rom[11897] = 16'hffff;
  rom[11898] = 16'hffff;
  rom[11899] = 16'hffff;
  rom[11900] = 16'hffff;
  rom[11901] = 16'hffff;
  rom[11902] = 16'hffff;
  rom[11903] = 16'hffff;
  rom[11904] = 16'hffff;
  rom[11905] = 16'hffff;
  rom[11906] = 16'hffff;
  rom[11907] = 16'hffff;
  rom[11908] = 16'hffff;
  rom[11909] = 16'hffff;
  rom[11910] = 16'hffff;
  rom[11911] = 16'hffff;
  rom[11912] = 16'hffff;
  rom[11913] = 16'hffff;
  rom[11914] = 16'hffff;
  rom[11915] = 16'hffff;
  rom[11916] = 16'hffff;
  rom[11917] = 16'hffff;
  rom[11918] = 16'hffff;
  rom[11919] = 16'hffff;
  rom[11920] = 16'hffff;
  rom[11921] = 16'hffff;
  rom[11922] = 16'hffff;
  rom[11923] = 16'hffff;
  rom[11924] = 16'hffff;
  rom[11925] = 16'hffff;
  rom[11926] = 16'hffff;
  rom[11927] = 16'hffff;
  rom[11928] = 16'hffff;
  rom[11929] = 16'hffff;
  rom[11930] = 16'hffff;
  rom[11931] = 16'hffff;
  rom[11932] = 16'hffff;
  rom[11933] = 16'hffff;
  rom[11934] = 16'hff9d;
  rom[11935] = 16'hac8e;
  rom[11936] = 16'h8326;
  rom[11937] = 16'hcd0c;
  rom[11938] = 16'hf5cc;
  rom[11939] = 16'hf5a9;
  rom[11940] = 16'hfda9;
  rom[11941] = 16'hfda8;
  rom[11942] = 16'hfd89;
  rom[11943] = 16'hf568;
  rom[11944] = 16'hfd88;
  rom[11945] = 16'hf567;
  rom[11946] = 16'hf548;
  rom[11947] = 16'hfd48;
  rom[11948] = 16'hfd49;
  rom[11949] = 16'hed6b;
  rom[11950] = 16'hb408;
  rom[11951] = 16'h7221;
  rom[11952] = 16'hc449;
  rom[11953] = 16'hcccd;
  rom[11954] = 16'h9bac;
  rom[11955] = 16'hff5d;
  rom[11956] = 16'hffff;
  rom[11957] = 16'hffff;
  rom[11958] = 16'hffff;
  rom[11959] = 16'hffff;
  rom[11960] = 16'hffff;
  rom[11961] = 16'hffff;
  rom[11962] = 16'hffff;
  rom[11963] = 16'hffff;
  rom[11964] = 16'hffff;
  rom[11965] = 16'hffff;
  rom[11966] = 16'hffff;
  rom[11967] = 16'hffff;
  rom[11968] = 16'hffff;
  rom[11969] = 16'hffff;
  rom[11970] = 16'hffff;
  rom[11971] = 16'hffff;
  rom[11972] = 16'hffff;
  rom[11973] = 16'hffff;
  rom[11974] = 16'hffff;
  rom[11975] = 16'hffff;
  rom[11976] = 16'hffff;
  rom[11977] = 16'hffff;
  rom[11978] = 16'hffff;
  rom[11979] = 16'hffff;
  rom[11980] = 16'hffff;
  rom[11981] = 16'hffff;
  rom[11982] = 16'hffff;
  rom[11983] = 16'hffff;
  rom[11984] = 16'hffff;
  rom[11985] = 16'hffff;
  rom[11986] = 16'hffff;
  rom[11987] = 16'hffff;
  rom[11988] = 16'hffff;
  rom[11989] = 16'hffff;
  rom[11990] = 16'hffff;
  rom[11991] = 16'hffff;
  rom[11992] = 16'hffff;
  rom[11993] = 16'hffff;
  rom[11994] = 16'hffff;
  rom[11995] = 16'hffff;
  rom[11996] = 16'hffff;
  rom[11997] = 16'hffff;
  rom[11998] = 16'hffff;
  rom[11999] = 16'hffff;
  rom[12000] = 16'hffff;
  rom[12001] = 16'hffff;
  rom[12002] = 16'hffff;
  rom[12003] = 16'hffff;
  rom[12004] = 16'hffff;
  rom[12005] = 16'hffff;
  rom[12006] = 16'hffff;
  rom[12007] = 16'hffff;
  rom[12008] = 16'hffff;
  rom[12009] = 16'hffff;
  rom[12010] = 16'hffff;
  rom[12011] = 16'hffff;
  rom[12012] = 16'hffff;
  rom[12013] = 16'hffff;
  rom[12014] = 16'hffff;
  rom[12015] = 16'hffff;
  rom[12016] = 16'hffff;
  rom[12017] = 16'hffff;
  rom[12018] = 16'hffff;
  rom[12019] = 16'hffff;
  rom[12020] = 16'hffff;
  rom[12021] = 16'hffff;
  rom[12022] = 16'hffff;
  rom[12023] = 16'hffff;
  rom[12024] = 16'hffff;
  rom[12025] = 16'hffff;
  rom[12026] = 16'hffff;
  rom[12027] = 16'hffff;
  rom[12028] = 16'hffff;
  rom[12029] = 16'hffff;
  rom[12030] = 16'hffff;
  rom[12031] = 16'hffff;
  rom[12032] = 16'hffff;
  rom[12033] = 16'hffff;
  rom[12034] = 16'hffff;
  rom[12035] = 16'hffff;
  rom[12036] = 16'hffff;
  rom[12037] = 16'hffdf;
  rom[12038] = 16'hfffe;
  rom[12039] = 16'h6ac8;
  rom[12040] = 16'h7b29;
  rom[12041] = 16'h72e8;
  rom[12042] = 16'h8bab;
  rom[12043] = 16'h7ae6;
  rom[12044] = 16'habe6;
  rom[12045] = 16'hf56a;
  rom[12046] = 16'hf507;
  rom[12047] = 16'hf548;
  rom[12048] = 16'hf568;
  rom[12049] = 16'hf568;
  rom[12050] = 16'hfd69;
  rom[12051] = 16'hfd68;
  rom[12052] = 16'hfd47;
  rom[12053] = 16'hfd69;
  rom[12054] = 16'hed48;
  rom[12055] = 16'hf5ab;
  rom[12056] = 16'hc4ca;
  rom[12057] = 16'h72e8;
  rom[12058] = 16'hc574;
  rom[12059] = 16'hfffe;
  rom[12060] = 16'hf79e;
  rom[12061] = 16'hffff;
  rom[12062] = 16'hffff;
  rom[12063] = 16'hffff;
  rom[12064] = 16'hffff;
  rom[12065] = 16'hffff;
  rom[12066] = 16'hffff;
  rom[12067] = 16'hffff;
  rom[12068] = 16'hffff;
  rom[12069] = 16'hffff;
  rom[12070] = 16'hffff;
  rom[12071] = 16'hffff;
  rom[12072] = 16'hffff;
  rom[12073] = 16'hffff;
  rom[12074] = 16'hffff;
  rom[12075] = 16'hffff;
  rom[12076] = 16'hffff;
  rom[12077] = 16'hffff;
  rom[12078] = 16'hffff;
  rom[12079] = 16'hffff;
  rom[12080] = 16'hffff;
  rom[12081] = 16'hffff;
  rom[12082] = 16'hffff;
  rom[12083] = 16'hffff;
  rom[12084] = 16'hffff;
  rom[12085] = 16'hffff;
  rom[12086] = 16'hffff;
  rom[12087] = 16'hffff;
  rom[12088] = 16'hffff;
  rom[12089] = 16'hffff;
  rom[12090] = 16'hffff;
  rom[12091] = 16'hffff;
  rom[12092] = 16'hffff;
  rom[12093] = 16'hffff;
  rom[12094] = 16'hffff;
  rom[12095] = 16'hffff;
  rom[12096] = 16'hffff;
  rom[12097] = 16'hffff;
  rom[12098] = 16'hffff;
  rom[12099] = 16'hffff;
  rom[12100] = 16'hffff;
  rom[12101] = 16'hffff;
  rom[12102] = 16'hffff;
  rom[12103] = 16'hffff;
  rom[12104] = 16'hffff;
  rom[12105] = 16'hffff;
  rom[12106] = 16'hffff;
  rom[12107] = 16'hffff;
  rom[12108] = 16'hffff;
  rom[12109] = 16'hffff;
  rom[12110] = 16'hffff;
  rom[12111] = 16'hffff;
  rom[12112] = 16'hffff;
  rom[12113] = 16'hffff;
  rom[12114] = 16'hffff;
  rom[12115] = 16'hffff;
  rom[12116] = 16'hffff;
  rom[12117] = 16'hffff;
  rom[12118] = 16'hffff;
  rom[12119] = 16'hffff;
  rom[12120] = 16'hffff;
  rom[12121] = 16'hffff;
  rom[12122] = 16'hffff;
  rom[12123] = 16'hffff;
  rom[12124] = 16'hffff;
  rom[12125] = 16'hffff;
  rom[12126] = 16'hffff;
  rom[12127] = 16'hffff;
  rom[12128] = 16'hffff;
  rom[12129] = 16'hffff;
  rom[12130] = 16'hffff;
  rom[12131] = 16'hffff;
  rom[12132] = 16'hffff;
  rom[12133] = 16'hffff;
  rom[12134] = 16'hffdf;
  rom[12135] = 16'hf75c;
  rom[12136] = 16'h942c;
  rom[12137] = 16'h9bc9;
  rom[12138] = 16'he5ce;
  rom[12139] = 16'he549;
  rom[12140] = 16'hf5a8;
  rom[12141] = 16'hfd68;
  rom[12142] = 16'hfd67;
  rom[12143] = 16'hfd87;
  rom[12144] = 16'hf567;
  rom[12145] = 16'hf587;
  rom[12146] = 16'hf568;
  rom[12147] = 16'hf549;
  rom[12148] = 16'hf528;
  rom[12149] = 16'hf549;
  rom[12150] = 16'hdcc9;
  rom[12151] = 16'ha345;
  rom[12152] = 16'hd4c8;
  rom[12153] = 16'hd50d;
  rom[12154] = 16'h93ac;
  rom[12155] = 16'hf73c;
  rom[12156] = 16'hffff;
  rom[12157] = 16'hffff;
  rom[12158] = 16'hffff;
  rom[12159] = 16'hffff;
  rom[12160] = 16'hffff;
  rom[12161] = 16'hffff;
  rom[12162] = 16'hffff;
  rom[12163] = 16'hffff;
  rom[12164] = 16'hffff;
  rom[12165] = 16'hffff;
  rom[12166] = 16'hffff;
  rom[12167] = 16'hffff;
  rom[12168] = 16'hffff;
  rom[12169] = 16'hffff;
  rom[12170] = 16'hffff;
  rom[12171] = 16'hffff;
  rom[12172] = 16'hffff;
  rom[12173] = 16'hffff;
  rom[12174] = 16'hffff;
  rom[12175] = 16'hffff;
  rom[12176] = 16'hffff;
  rom[12177] = 16'hffff;
  rom[12178] = 16'hffff;
  rom[12179] = 16'hffff;
  rom[12180] = 16'hffff;
  rom[12181] = 16'hffff;
  rom[12182] = 16'hffff;
  rom[12183] = 16'hffff;
  rom[12184] = 16'hffff;
  rom[12185] = 16'hffff;
  rom[12186] = 16'hffff;
  rom[12187] = 16'hffff;
  rom[12188] = 16'hffff;
  rom[12189] = 16'hffff;
  rom[12190] = 16'hffff;
  rom[12191] = 16'hffff;
  rom[12192] = 16'hffff;
  rom[12193] = 16'hffff;
  rom[12194] = 16'hffff;
  rom[12195] = 16'hffff;
  rom[12196] = 16'hffff;
  rom[12197] = 16'hffff;
  rom[12198] = 16'hffff;
  rom[12199] = 16'hffff;
  rom[12200] = 16'hffff;
  rom[12201] = 16'hffff;
  rom[12202] = 16'hffff;
  rom[12203] = 16'hffff;
  rom[12204] = 16'hffff;
  rom[12205] = 16'hffff;
  rom[12206] = 16'hffff;
  rom[12207] = 16'hffff;
  rom[12208] = 16'hffff;
  rom[12209] = 16'hffff;
  rom[12210] = 16'hffff;
  rom[12211] = 16'hffff;
  rom[12212] = 16'hffff;
  rom[12213] = 16'hffff;
  rom[12214] = 16'hffff;
  rom[12215] = 16'hffff;
  rom[12216] = 16'hffff;
  rom[12217] = 16'hffff;
  rom[12218] = 16'hffff;
  rom[12219] = 16'hffff;
  rom[12220] = 16'hffff;
  rom[12221] = 16'hffff;
  rom[12222] = 16'hffff;
  rom[12223] = 16'hffff;
  rom[12224] = 16'hffff;
  rom[12225] = 16'hffff;
  rom[12226] = 16'hffff;
  rom[12227] = 16'hffff;
  rom[12228] = 16'hffff;
  rom[12229] = 16'hffff;
  rom[12230] = 16'hffff;
  rom[12231] = 16'hffff;
  rom[12232] = 16'hffff;
  rom[12233] = 16'hffff;
  rom[12234] = 16'hffff;
  rom[12235] = 16'hffff;
  rom[12236] = 16'hffff;
  rom[12237] = 16'hffff;
  rom[12238] = 16'hffde;
  rom[12239] = 16'ha46e;
  rom[12240] = 16'ha42c;
  rom[12241] = 16'hc4ef;
  rom[12242] = 16'habea;
  rom[12243] = 16'h9ba6;
  rom[12244] = 16'hcca8;
  rom[12245] = 16'hfd6a;
  rom[12246] = 16'hfd69;
  rom[12247] = 16'hf568;
  rom[12248] = 16'hfd68;
  rom[12249] = 16'hf568;
  rom[12250] = 16'hfd68;
  rom[12251] = 16'hfd68;
  rom[12252] = 16'hfd89;
  rom[12253] = 16'hf528;
  rom[12254] = 16'hf58b;
  rom[12255] = 16'hdd6c;
  rom[12256] = 16'h8b88;
  rom[12257] = 16'hacf1;
  rom[12258] = 16'hffbd;
  rom[12259] = 16'hffff;
  rom[12260] = 16'hffdf;
  rom[12261] = 16'hffff;
  rom[12262] = 16'hffff;
  rom[12263] = 16'hffff;
  rom[12264] = 16'hffff;
  rom[12265] = 16'hffff;
  rom[12266] = 16'hffff;
  rom[12267] = 16'hffff;
  rom[12268] = 16'hffff;
  rom[12269] = 16'hffff;
  rom[12270] = 16'hffff;
  rom[12271] = 16'hffff;
  rom[12272] = 16'hffff;
  rom[12273] = 16'hffff;
  rom[12274] = 16'hffff;
  rom[12275] = 16'hffff;
  rom[12276] = 16'hffff;
  rom[12277] = 16'hffff;
  rom[12278] = 16'hffff;
  rom[12279] = 16'hffff;
  rom[12280] = 16'hffff;
  rom[12281] = 16'hffff;
  rom[12282] = 16'hffff;
  rom[12283] = 16'hffff;
  rom[12284] = 16'hffff;
  rom[12285] = 16'hffff;
  rom[12286] = 16'hffff;
  rom[12287] = 16'hffff;
  rom[12288] = 16'hffff;
  rom[12289] = 16'hffff;
  rom[12290] = 16'hffff;
  rom[12291] = 16'hffff;
  rom[12292] = 16'hffff;
  rom[12293] = 16'hffff;
  rom[12294] = 16'hffff;
  rom[12295] = 16'hffff;
  rom[12296] = 16'hffff;
  rom[12297] = 16'hffff;
  rom[12298] = 16'hffff;
  rom[12299] = 16'hffff;
  rom[12300] = 16'hffff;
  rom[12301] = 16'hffff;
  rom[12302] = 16'hffff;
  rom[12303] = 16'hffff;
  rom[12304] = 16'hffff;
  rom[12305] = 16'hffff;
  rom[12306] = 16'hffff;
  rom[12307] = 16'hffff;
  rom[12308] = 16'hffff;
  rom[12309] = 16'hffff;
  rom[12310] = 16'hffff;
  rom[12311] = 16'hffff;
  rom[12312] = 16'hffff;
  rom[12313] = 16'hffff;
  rom[12314] = 16'hffff;
  rom[12315] = 16'hffff;
  rom[12316] = 16'hffff;
  rom[12317] = 16'hffff;
  rom[12318] = 16'hffff;
  rom[12319] = 16'hffff;
  rom[12320] = 16'hffff;
  rom[12321] = 16'hffff;
  rom[12322] = 16'hffff;
  rom[12323] = 16'hffff;
  rom[12324] = 16'hffff;
  rom[12325] = 16'hffff;
  rom[12326] = 16'hffff;
  rom[12327] = 16'hffff;
  rom[12328] = 16'hffff;
  rom[12329] = 16'hffff;
  rom[12330] = 16'hffff;
  rom[12331] = 16'hffff;
  rom[12332] = 16'hffff;
  rom[12333] = 16'hffff;
  rom[12334] = 16'hffff;
  rom[12335] = 16'hffff;
  rom[12336] = 16'he6d9;
  rom[12337] = 16'h8369;
  rom[12338] = 16'hbcab;
  rom[12339] = 16'hedcd;
  rom[12340] = 16'hf58a;
  rom[12341] = 16'hf568;
  rom[12342] = 16'hfd68;
  rom[12343] = 16'hfd67;
  rom[12344] = 16'hfd67;
  rom[12345] = 16'hf567;
  rom[12346] = 16'hf569;
  rom[12347] = 16'hf549;
  rom[12348] = 16'hfd6a;
  rom[12349] = 16'hf548;
  rom[12350] = 16'hfd6a;
  rom[12351] = 16'hdcc9;
  rom[12352] = 16'hed6a;
  rom[12353] = 16'hdd4b;
  rom[12354] = 16'h936b;
  rom[12355] = 16'hde79;
  rom[12356] = 16'hffff;
  rom[12357] = 16'hffff;
  rom[12358] = 16'hffff;
  rom[12359] = 16'hffff;
  rom[12360] = 16'hffff;
  rom[12361] = 16'hffff;
  rom[12362] = 16'hffff;
  rom[12363] = 16'hffff;
  rom[12364] = 16'hffff;
  rom[12365] = 16'hffff;
  rom[12366] = 16'hffff;
  rom[12367] = 16'hffff;
  rom[12368] = 16'hffff;
  rom[12369] = 16'hffff;
  rom[12370] = 16'hffff;
  rom[12371] = 16'hffff;
  rom[12372] = 16'hffff;
  rom[12373] = 16'hffff;
  rom[12374] = 16'hffff;
  rom[12375] = 16'hffff;
  rom[12376] = 16'hffff;
  rom[12377] = 16'hffff;
  rom[12378] = 16'hffff;
  rom[12379] = 16'hffff;
  rom[12380] = 16'hffff;
  rom[12381] = 16'hffff;
  rom[12382] = 16'hffff;
  rom[12383] = 16'hffff;
  rom[12384] = 16'hffff;
  rom[12385] = 16'hffff;
  rom[12386] = 16'hffff;
  rom[12387] = 16'hffff;
  rom[12388] = 16'hffff;
  rom[12389] = 16'hffff;
  rom[12390] = 16'hffff;
  rom[12391] = 16'hffff;
  rom[12392] = 16'hffff;
  rom[12393] = 16'hffff;
  rom[12394] = 16'hffff;
  rom[12395] = 16'hffff;
  rom[12396] = 16'hffff;
  rom[12397] = 16'hffff;
  rom[12398] = 16'hffff;
  rom[12399] = 16'hffff;
  rom[12400] = 16'hffff;
  rom[12401] = 16'hffff;
  rom[12402] = 16'hffff;
  rom[12403] = 16'hffff;
  rom[12404] = 16'hffff;
  rom[12405] = 16'hffff;
  rom[12406] = 16'hffff;
  rom[12407] = 16'hffff;
  rom[12408] = 16'hffff;
  rom[12409] = 16'hffff;
  rom[12410] = 16'hffff;
  rom[12411] = 16'hffff;
  rom[12412] = 16'hffff;
  rom[12413] = 16'hffff;
  rom[12414] = 16'hffff;
  rom[12415] = 16'hffff;
  rom[12416] = 16'hffff;
  rom[12417] = 16'hffff;
  rom[12418] = 16'hffff;
  rom[12419] = 16'hffff;
  rom[12420] = 16'hffff;
  rom[12421] = 16'hffff;
  rom[12422] = 16'hffff;
  rom[12423] = 16'hffff;
  rom[12424] = 16'hffff;
  rom[12425] = 16'hffff;
  rom[12426] = 16'hffff;
  rom[12427] = 16'hffff;
  rom[12428] = 16'hffff;
  rom[12429] = 16'hffff;
  rom[12430] = 16'hffff;
  rom[12431] = 16'hffff;
  rom[12432] = 16'hffff;
  rom[12433] = 16'hffff;
  rom[12434] = 16'hffff;
  rom[12435] = 16'hffff;
  rom[12436] = 16'hffdf;
  rom[12437] = 16'hffff;
  rom[12438] = 16'hffde;
  rom[12439] = 16'hd5f5;
  rom[12440] = 16'h82c6;
  rom[12441] = 16'hd52e;
  rom[12442] = 16'he58d;
  rom[12443] = 16'hedac;
  rom[12444] = 16'hfd8a;
  rom[12445] = 16'hecc9;
  rom[12446] = 16'hf529;
  rom[12447] = 16'hf549;
  rom[12448] = 16'hf568;
  rom[12449] = 16'hf588;
  rom[12450] = 16'hf567;
  rom[12451] = 16'hfd47;
  rom[12452] = 16'hfd28;
  rom[12453] = 16'hfd8c;
  rom[12454] = 16'he56c;
  rom[12455] = 16'hbccc;
  rom[12456] = 16'h8389;
  rom[12457] = 16'hf77c;
  rom[12458] = 16'hffde;
  rom[12459] = 16'hffff;
  rom[12460] = 16'hffff;
  rom[12461] = 16'hffff;
  rom[12462] = 16'hffff;
  rom[12463] = 16'hffff;
  rom[12464] = 16'hffff;
  rom[12465] = 16'hffff;
  rom[12466] = 16'hffff;
  rom[12467] = 16'hffff;
  rom[12468] = 16'hffff;
  rom[12469] = 16'hffff;
  rom[12470] = 16'hffff;
  rom[12471] = 16'hffff;
  rom[12472] = 16'hffff;
  rom[12473] = 16'hffff;
  rom[12474] = 16'hffff;
  rom[12475] = 16'hffff;
  rom[12476] = 16'hffff;
  rom[12477] = 16'hffff;
  rom[12478] = 16'hffff;
  rom[12479] = 16'hffff;
  rom[12480] = 16'hffff;
  rom[12481] = 16'hffff;
  rom[12482] = 16'hffff;
  rom[12483] = 16'hffff;
  rom[12484] = 16'hffff;
  rom[12485] = 16'hffff;
  rom[12486] = 16'hffff;
  rom[12487] = 16'hffff;
  rom[12488] = 16'hffff;
  rom[12489] = 16'hffff;
  rom[12490] = 16'hffff;
  rom[12491] = 16'hffff;
  rom[12492] = 16'hffff;
  rom[12493] = 16'hffff;
  rom[12494] = 16'hffff;
  rom[12495] = 16'hffff;
  rom[12496] = 16'hffff;
  rom[12497] = 16'hffff;
  rom[12498] = 16'hffff;
  rom[12499] = 16'hffff;
  rom[12500] = 16'hffff;
  rom[12501] = 16'hffff;
  rom[12502] = 16'hffff;
  rom[12503] = 16'hffff;
  rom[12504] = 16'hffff;
  rom[12505] = 16'hffff;
  rom[12506] = 16'hffff;
  rom[12507] = 16'hffff;
  rom[12508] = 16'hffdf;
  rom[12509] = 16'hffff;
  rom[12510] = 16'hffff;
  rom[12511] = 16'hffff;
  rom[12512] = 16'hffff;
  rom[12513] = 16'hffff;
  rom[12514] = 16'hffff;
  rom[12515] = 16'hffff;
  rom[12516] = 16'hffff;
  rom[12517] = 16'hffff;
  rom[12518] = 16'hffff;
  rom[12519] = 16'hffff;
  rom[12520] = 16'hffff;
  rom[12521] = 16'hffff;
  rom[12522] = 16'hffff;
  rom[12523] = 16'hffff;
  rom[12524] = 16'hffff;
  rom[12525] = 16'hffff;
  rom[12526] = 16'hffff;
  rom[12527] = 16'hffff;
  rom[12528] = 16'hffff;
  rom[12529] = 16'hffff;
  rom[12530] = 16'hffff;
  rom[12531] = 16'hffff;
  rom[12532] = 16'hffff;
  rom[12533] = 16'hffff;
  rom[12534] = 16'hffff;
  rom[12535] = 16'hffff;
  rom[12536] = 16'hffde;
  rom[12537] = 16'hbd93;
  rom[12538] = 16'h72e6;
  rom[12539] = 16'hcd0c;
  rom[12540] = 16'hed8b;
  rom[12541] = 16'hfd69;
  rom[12542] = 16'hfd67;
  rom[12543] = 16'hfd67;
  rom[12544] = 16'hfd67;
  rom[12545] = 16'hfd88;
  rom[12546] = 16'hed48;
  rom[12547] = 16'hfd6a;
  rom[12548] = 16'hf528;
  rom[12549] = 16'hf506;
  rom[12550] = 16'hf568;
  rom[12551] = 16'hfd6a;
  rom[12552] = 16'hed68;
  rom[12553] = 16'hdd4b;
  rom[12554] = 16'h7ac6;
  rom[12555] = 16'hd657;
  rom[12556] = 16'hffff;
  rom[12557] = 16'hffff;
  rom[12558] = 16'hffff;
  rom[12559] = 16'hffff;
  rom[12560] = 16'hffff;
  rom[12561] = 16'hffff;
  rom[12562] = 16'hffff;
  rom[12563] = 16'hffff;
  rom[12564] = 16'hffff;
  rom[12565] = 16'hffff;
  rom[12566] = 16'hffff;
  rom[12567] = 16'hffff;
  rom[12568] = 16'hffff;
  rom[12569] = 16'hffff;
  rom[12570] = 16'hffff;
  rom[12571] = 16'hffff;
  rom[12572] = 16'hffff;
  rom[12573] = 16'hffff;
  rom[12574] = 16'hffff;
  rom[12575] = 16'hffff;
  rom[12576] = 16'hffff;
  rom[12577] = 16'hffff;
  rom[12578] = 16'hffff;
  rom[12579] = 16'hffff;
  rom[12580] = 16'hffff;
  rom[12581] = 16'hffff;
  rom[12582] = 16'hffff;
  rom[12583] = 16'hffff;
  rom[12584] = 16'hffff;
  rom[12585] = 16'hffff;
  rom[12586] = 16'hffff;
  rom[12587] = 16'hffff;
  rom[12588] = 16'hffff;
  rom[12589] = 16'hffff;
  rom[12590] = 16'hffff;
  rom[12591] = 16'hffff;
  rom[12592] = 16'hffff;
  rom[12593] = 16'hffff;
  rom[12594] = 16'hffff;
  rom[12595] = 16'hffff;
  rom[12596] = 16'hffff;
  rom[12597] = 16'hffff;
  rom[12598] = 16'hffff;
  rom[12599] = 16'hffff;
  rom[12600] = 16'hffff;
  rom[12601] = 16'hffff;
  rom[12602] = 16'hffff;
  rom[12603] = 16'hffff;
  rom[12604] = 16'hffff;
  rom[12605] = 16'hffff;
  rom[12606] = 16'hffff;
  rom[12607] = 16'hffff;
  rom[12608] = 16'hffff;
  rom[12609] = 16'hffff;
  rom[12610] = 16'hffff;
  rom[12611] = 16'hffff;
  rom[12612] = 16'hffff;
  rom[12613] = 16'hffff;
  rom[12614] = 16'hffff;
  rom[12615] = 16'hffff;
  rom[12616] = 16'hffff;
  rom[12617] = 16'hffff;
  rom[12618] = 16'hffff;
  rom[12619] = 16'hffff;
  rom[12620] = 16'hffff;
  rom[12621] = 16'hffff;
  rom[12622] = 16'hffff;
  rom[12623] = 16'hffff;
  rom[12624] = 16'hffff;
  rom[12625] = 16'hffff;
  rom[12626] = 16'hffff;
  rom[12627] = 16'hffff;
  rom[12628] = 16'hffff;
  rom[12629] = 16'hffff;
  rom[12630] = 16'hffff;
  rom[12631] = 16'hffff;
  rom[12632] = 16'hffff;
  rom[12633] = 16'hffff;
  rom[12634] = 16'hffff;
  rom[12635] = 16'hffff;
  rom[12636] = 16'hffff;
  rom[12637] = 16'hffff;
  rom[12638] = 16'hffff;
  rom[12639] = 16'hf6da;
  rom[12640] = 16'h82e8;
  rom[12641] = 16'hbc4b;
  rom[12642] = 16'he58d;
  rom[12643] = 16'hed6a;
  rom[12644] = 16'hfd2a;
  rom[12645] = 16'hfd29;
  rom[12646] = 16'hfd6a;
  rom[12647] = 16'hf549;
  rom[12648] = 16'hf589;
  rom[12649] = 16'hf566;
  rom[12650] = 16'hfd86;
  rom[12651] = 16'hfd67;
  rom[12652] = 16'hfd69;
  rom[12653] = 16'hf58c;
  rom[12654] = 16'hd50e;
  rom[12655] = 16'h8308;
  rom[12656] = 16'hcdd5;
  rom[12657] = 16'hffff;
  rom[12658] = 16'hffff;
  rom[12659] = 16'hffff;
  rom[12660] = 16'hffff;
  rom[12661] = 16'hffff;
  rom[12662] = 16'hffff;
  rom[12663] = 16'hffff;
  rom[12664] = 16'hffff;
  rom[12665] = 16'hffff;
  rom[12666] = 16'hffff;
  rom[12667] = 16'hffff;
  rom[12668] = 16'hffff;
  rom[12669] = 16'hffff;
  rom[12670] = 16'hffff;
  rom[12671] = 16'hffff;
  rom[12672] = 16'hffff;
  rom[12673] = 16'hffff;
  rom[12674] = 16'hffff;
  rom[12675] = 16'hffff;
  rom[12676] = 16'hffff;
  rom[12677] = 16'hffff;
  rom[12678] = 16'hffff;
  rom[12679] = 16'hffff;
  rom[12680] = 16'hffff;
  rom[12681] = 16'hffff;
  rom[12682] = 16'hffff;
  rom[12683] = 16'hffff;
  rom[12684] = 16'hffff;
  rom[12685] = 16'hffff;
  rom[12686] = 16'hffff;
  rom[12687] = 16'hffff;
  rom[12688] = 16'hffff;
  rom[12689] = 16'hffff;
  rom[12690] = 16'hffff;
  rom[12691] = 16'hffff;
  rom[12692] = 16'hffff;
  rom[12693] = 16'hffff;
  rom[12694] = 16'hffff;
  rom[12695] = 16'hffff;
  rom[12696] = 16'hffff;
  rom[12697] = 16'hffff;
  rom[12698] = 16'hffff;
  rom[12699] = 16'hffff;
  rom[12700] = 16'hffff;
  rom[12701] = 16'hffff;
  rom[12702] = 16'hffff;
  rom[12703] = 16'hffff;
  rom[12704] = 16'hffff;
  rom[12705] = 16'hffff;
  rom[12706] = 16'hffff;
  rom[12707] = 16'hffff;
  rom[12708] = 16'hffff;
  rom[12709] = 16'hffff;
  rom[12710] = 16'hffff;
  rom[12711] = 16'hffff;
  rom[12712] = 16'hffff;
  rom[12713] = 16'hffff;
  rom[12714] = 16'hffff;
  rom[12715] = 16'hffff;
  rom[12716] = 16'hffff;
  rom[12717] = 16'hffff;
  rom[12718] = 16'hffff;
  rom[12719] = 16'hffff;
  rom[12720] = 16'hffff;
  rom[12721] = 16'hffff;
  rom[12722] = 16'hffff;
  rom[12723] = 16'hffff;
  rom[12724] = 16'hffff;
  rom[12725] = 16'hffff;
  rom[12726] = 16'hffff;
  rom[12727] = 16'hffff;
  rom[12728] = 16'hffff;
  rom[12729] = 16'hffff;
  rom[12730] = 16'hffff;
  rom[12731] = 16'hffff;
  rom[12732] = 16'hffff;
  rom[12733] = 16'hffff;
  rom[12734] = 16'hffff;
  rom[12735] = 16'hffff;
  rom[12736] = 16'hffff;
  rom[12737] = 16'hf77c;
  rom[12738] = 16'h8bcb;
  rom[12739] = 16'ha3e9;
  rom[12740] = 16'hed8d;
  rom[12741] = 16'hf58b;
  rom[12742] = 16'hfd68;
  rom[12743] = 16'hfd47;
  rom[12744] = 16'hfd68;
  rom[12745] = 16'hfd48;
  rom[12746] = 16'hf569;
  rom[12747] = 16'hf549;
  rom[12748] = 16'hfd49;
  rom[12749] = 16'hfd67;
  rom[12750] = 16'hfd47;
  rom[12751] = 16'hf528;
  rom[12752] = 16'hf569;
  rom[12753] = 16'he52a;
  rom[12754] = 16'h82e7;
  rom[12755] = 16'hcdf6;
  rom[12756] = 16'hffff;
  rom[12757] = 16'hffff;
  rom[12758] = 16'hffff;
  rom[12759] = 16'hffff;
  rom[12760] = 16'hffff;
  rom[12761] = 16'hffff;
  rom[12762] = 16'hffff;
  rom[12763] = 16'hffff;
  rom[12764] = 16'hffff;
  rom[12765] = 16'hffff;
  rom[12766] = 16'hffff;
  rom[12767] = 16'hffff;
  rom[12768] = 16'hffff;
  rom[12769] = 16'hffff;
  rom[12770] = 16'hffff;
  rom[12771] = 16'hffff;
  rom[12772] = 16'hffff;
  rom[12773] = 16'hffff;
  rom[12774] = 16'hffff;
  rom[12775] = 16'hffff;
  rom[12776] = 16'hffff;
  rom[12777] = 16'hffff;
  rom[12778] = 16'hffff;
  rom[12779] = 16'hffff;
  rom[12780] = 16'hffff;
  rom[12781] = 16'hffff;
  rom[12782] = 16'hffff;
  rom[12783] = 16'hffff;
  rom[12784] = 16'hffff;
  rom[12785] = 16'hffff;
  rom[12786] = 16'hffff;
  rom[12787] = 16'hffff;
  rom[12788] = 16'hffff;
  rom[12789] = 16'hffff;
  rom[12790] = 16'hffff;
  rom[12791] = 16'hffff;
  rom[12792] = 16'hffff;
  rom[12793] = 16'hffff;
  rom[12794] = 16'hffff;
  rom[12795] = 16'hffff;
  rom[12796] = 16'hffff;
  rom[12797] = 16'hffff;
  rom[12798] = 16'hffff;
  rom[12799] = 16'hffff;
  rom[12800] = 16'hffff;
  rom[12801] = 16'hffff;
  rom[12802] = 16'hffff;
  rom[12803] = 16'hffff;
  rom[12804] = 16'hffff;
  rom[12805] = 16'hffff;
  rom[12806] = 16'hffff;
  rom[12807] = 16'hffff;
  rom[12808] = 16'hffff;
  rom[12809] = 16'hffff;
  rom[12810] = 16'hffff;
  rom[12811] = 16'hffff;
  rom[12812] = 16'hffff;
  rom[12813] = 16'hffff;
  rom[12814] = 16'hffff;
  rom[12815] = 16'hffff;
  rom[12816] = 16'hffff;
  rom[12817] = 16'hffff;
  rom[12818] = 16'hffff;
  rom[12819] = 16'hffff;
  rom[12820] = 16'hffff;
  rom[12821] = 16'hffff;
  rom[12822] = 16'hffff;
  rom[12823] = 16'hffff;
  rom[12824] = 16'hffff;
  rom[12825] = 16'hffff;
  rom[12826] = 16'hffff;
  rom[12827] = 16'hffff;
  rom[12828] = 16'hffff;
  rom[12829] = 16'hffff;
  rom[12830] = 16'hffff;
  rom[12831] = 16'hffff;
  rom[12832] = 16'hffff;
  rom[12833] = 16'hffff;
  rom[12834] = 16'hffff;
  rom[12835] = 16'hffff;
  rom[12836] = 16'hfffe;
  rom[12837] = 16'hffff;
  rom[12838] = 16'hffdf;
  rom[12839] = 16'hff9e;
  rom[12840] = 16'hcd32;
  rom[12841] = 16'h7263;
  rom[12842] = 16'hdd6c;
  rom[12843] = 16'hdd09;
  rom[12844] = 16'hf528;
  rom[12845] = 16'hfd29;
  rom[12846] = 16'hf508;
  rom[12847] = 16'hf569;
  rom[12848] = 16'hed69;
  rom[12849] = 16'hfd88;
  rom[12850] = 16'hfd46;
  rom[12851] = 16'hfd67;
  rom[12852] = 16'hf58a;
  rom[12853] = 16'he56d;
  rom[12854] = 16'h9bca;
  rom[12855] = 16'h8b8c;
  rom[12856] = 16'hff9d;
  rom[12857] = 16'hffff;
  rom[12858] = 16'hffff;
  rom[12859] = 16'hffff;
  rom[12860] = 16'hffff;
  rom[12861] = 16'hffff;
  rom[12862] = 16'hffff;
  rom[12863] = 16'hffff;
  rom[12864] = 16'hffff;
  rom[12865] = 16'hffff;
  rom[12866] = 16'hffff;
  rom[12867] = 16'hffff;
  rom[12868] = 16'hffff;
  rom[12869] = 16'hffff;
  rom[12870] = 16'hffff;
  rom[12871] = 16'hffff;
  rom[12872] = 16'hffff;
  rom[12873] = 16'hffff;
  rom[12874] = 16'hffff;
  rom[12875] = 16'hffff;
  rom[12876] = 16'hffff;
  rom[12877] = 16'hffff;
  rom[12878] = 16'hffbf;
  rom[12879] = 16'hffff;
  rom[12880] = 16'hffdf;
  rom[12881] = 16'hffff;
  rom[12882] = 16'hffff;
  rom[12883] = 16'hffff;
  rom[12884] = 16'hffff;
  rom[12885] = 16'hffff;
  rom[12886] = 16'hffff;
  rom[12887] = 16'hffff;
  rom[12888] = 16'hffff;
  rom[12889] = 16'hffff;
  rom[12890] = 16'hffff;
  rom[12891] = 16'hffff;
  rom[12892] = 16'hffff;
  rom[12893] = 16'hffff;
  rom[12894] = 16'hffff;
  rom[12895] = 16'hffff;
  rom[12896] = 16'hffff;
  rom[12897] = 16'hffff;
  rom[12898] = 16'hffff;
  rom[12899] = 16'hffff;
  rom[12900] = 16'hffff;
  rom[12901] = 16'hffff;
  rom[12902] = 16'hffff;
  rom[12903] = 16'hffff;
  rom[12904] = 16'hffff;
  rom[12905] = 16'hffff;
  rom[12906] = 16'hffff;
  rom[12907] = 16'hffff;
  rom[12908] = 16'hffff;
  rom[12909] = 16'hffff;
  rom[12910] = 16'hffff;
  rom[12911] = 16'hffff;
  rom[12912] = 16'hffdf;
  rom[12913] = 16'hffff;
  rom[12914] = 16'hffdf;
  rom[12915] = 16'hffff;
  rom[12916] = 16'hffff;
  rom[12917] = 16'hffff;
  rom[12918] = 16'hffdf;
  rom[12919] = 16'hffff;
  rom[12920] = 16'hffff;
  rom[12921] = 16'hffff;
  rom[12922] = 16'hffff;
  rom[12923] = 16'hffff;
  rom[12924] = 16'hffff;
  rom[12925] = 16'hffff;
  rom[12926] = 16'hffff;
  rom[12927] = 16'hffff;
  rom[12928] = 16'hffff;
  rom[12929] = 16'hffff;
  rom[12930] = 16'hffff;
  rom[12931] = 16'hffff;
  rom[12932] = 16'hfffe;
  rom[12933] = 16'hffff;
  rom[12934] = 16'hffff;
  rom[12935] = 16'hffff;
  rom[12936] = 16'hffff;
  rom[12937] = 16'hfffe;
  rom[12938] = 16'hde97;
  rom[12939] = 16'h8b8a;
  rom[12940] = 16'hcd2d;
  rom[12941] = 16'hed4a;
  rom[12942] = 16'hfd69;
  rom[12943] = 16'hfd68;
  rom[12944] = 16'hfd47;
  rom[12945] = 16'hfd69;
  rom[12946] = 16'hf549;
  rom[12947] = 16'hf568;
  rom[12948] = 16'hf528;
  rom[12949] = 16'hfd47;
  rom[12950] = 16'hf547;
  rom[12951] = 16'hf549;
  rom[12952] = 16'hed48;
  rom[12953] = 16'he54a;
  rom[12954] = 16'h82c6;
  rom[12955] = 16'hc595;
  rom[12956] = 16'hffdf;
  rom[12957] = 16'hffff;
  rom[12958] = 16'hffff;
  rom[12959] = 16'hffff;
  rom[12960] = 16'hffff;
  rom[12961] = 16'hffff;
  rom[12962] = 16'hffff;
  rom[12963] = 16'hffff;
  rom[12964] = 16'hffff;
  rom[12965] = 16'hffff;
  rom[12966] = 16'hffff;
  rom[12967] = 16'hffff;
  rom[12968] = 16'hffff;
  rom[12969] = 16'hffff;
  rom[12970] = 16'hffff;
  rom[12971] = 16'hffff;
  rom[12972] = 16'hffff;
  rom[12973] = 16'hffff;
  rom[12974] = 16'hffff;
  rom[12975] = 16'hffff;
  rom[12976] = 16'hffff;
  rom[12977] = 16'hffff;
  rom[12978] = 16'hffff;
  rom[12979] = 16'hffff;
  rom[12980] = 16'hffff;
  rom[12981] = 16'hffff;
  rom[12982] = 16'hffff;
  rom[12983] = 16'hffff;
  rom[12984] = 16'hffff;
  rom[12985] = 16'hffff;
  rom[12986] = 16'hffff;
  rom[12987] = 16'hffff;
  rom[12988] = 16'hffff;
  rom[12989] = 16'hffff;
  rom[12990] = 16'hffff;
  rom[12991] = 16'hffff;
  rom[12992] = 16'hffff;
  rom[12993] = 16'hffff;
  rom[12994] = 16'hffff;
  rom[12995] = 16'hffff;
  rom[12996] = 16'hffff;
  rom[12997] = 16'hffff;
  rom[12998] = 16'hffff;
  rom[12999] = 16'hffff;
  rom[13000] = 16'hffff;
  rom[13001] = 16'hffff;
  rom[13002] = 16'hffff;
  rom[13003] = 16'hffff;
  rom[13004] = 16'hffff;
  rom[13005] = 16'hffff;
  rom[13006] = 16'hffff;
  rom[13007] = 16'hffff;
  rom[13008] = 16'hffff;
  rom[13009] = 16'hffff;
  rom[13010] = 16'hffff;
  rom[13011] = 16'hffff;
  rom[13012] = 16'hffff;
  rom[13013] = 16'hffff;
  rom[13014] = 16'hffff;
  rom[13015] = 16'hffff;
  rom[13016] = 16'hffff;
  rom[13017] = 16'hffff;
  rom[13018] = 16'hffff;
  rom[13019] = 16'hffff;
  rom[13020] = 16'hffff;
  rom[13021] = 16'hffff;
  rom[13022] = 16'hffff;
  rom[13023] = 16'hffff;
  rom[13024] = 16'hffff;
  rom[13025] = 16'hffff;
  rom[13026] = 16'hffff;
  rom[13027] = 16'hffff;
  rom[13028] = 16'hffff;
  rom[13029] = 16'hffff;
  rom[13030] = 16'hffff;
  rom[13031] = 16'hffff;
  rom[13032] = 16'hffff;
  rom[13033] = 16'hffff;
  rom[13034] = 16'hffff;
  rom[13035] = 16'hffff;
  rom[13036] = 16'hffff;
  rom[13037] = 16'hffff;
  rom[13038] = 16'hffff;
  rom[13039] = 16'hffbf;
  rom[13040] = 16'hff1b;
  rom[13041] = 16'h9beb;
  rom[13042] = 16'h9386;
  rom[13043] = 16'hfdcc;
  rom[13044] = 16'hfd49;
  rom[13045] = 16'hfd48;
  rom[13046] = 16'hfd69;
  rom[13047] = 16'hf569;
  rom[13048] = 16'hf569;
  rom[13049] = 16'hf547;
  rom[13050] = 16'hfd47;
  rom[13051] = 16'hfd48;
  rom[13052] = 16'hfdcc;
  rom[13053] = 16'hcd0c;
  rom[13054] = 16'h8b6a;
  rom[13055] = 16'hde58;
  rom[13056] = 16'hffbf;
  rom[13057] = 16'hffff;
  rom[13058] = 16'hffff;
  rom[13059] = 16'hffff;
  rom[13060] = 16'hffff;
  rom[13061] = 16'hffff;
  rom[13062] = 16'hffff;
  rom[13063] = 16'hffff;
  rom[13064] = 16'hffff;
  rom[13065] = 16'hffff;
  rom[13066] = 16'hffff;
  rom[13067] = 16'hffff;
  rom[13068] = 16'hffff;
  rom[13069] = 16'hffff;
  rom[13070] = 16'hffff;
  rom[13071] = 16'hffff;
  rom[13072] = 16'hffff;
  rom[13073] = 16'hffff;
  rom[13074] = 16'hffff;
  rom[13075] = 16'hffff;
  rom[13076] = 16'hffff;
  rom[13077] = 16'hffff;
  rom[13078] = 16'hffff;
  rom[13079] = 16'hffff;
  rom[13080] = 16'hffff;
  rom[13081] = 16'hffff;
  rom[13082] = 16'hffff;
  rom[13083] = 16'hffff;
  rom[13084] = 16'hffff;
  rom[13085] = 16'hffff;
  rom[13086] = 16'hffff;
  rom[13087] = 16'hffff;
  rom[13088] = 16'hffff;
  rom[13089] = 16'hffff;
  rom[13090] = 16'hffff;
  rom[13091] = 16'hffff;
  rom[13092] = 16'hffff;
  rom[13093] = 16'hffff;
  rom[13094] = 16'hffff;
  rom[13095] = 16'hffff;
  rom[13096] = 16'hffff;
  rom[13097] = 16'hffff;
  rom[13098] = 16'hffff;
  rom[13099] = 16'hffff;
  rom[13100] = 16'hffff;
  rom[13101] = 16'hffff;
  rom[13102] = 16'hffff;
  rom[13103] = 16'hffff;
  rom[13104] = 16'hffff;
  rom[13105] = 16'hffff;
  rom[13106] = 16'hffff;
  rom[13107] = 16'hffff;
  rom[13108] = 16'hffff;
  rom[13109] = 16'hffdf;
  rom[13110] = 16'hffff;
  rom[13111] = 16'hffdf;
  rom[13112] = 16'hffff;
  rom[13113] = 16'hffff;
  rom[13114] = 16'hffff;
  rom[13115] = 16'hffff;
  rom[13116] = 16'hffff;
  rom[13117] = 16'hffff;
  rom[13118] = 16'hffff;
  rom[13119] = 16'hffff;
  rom[13120] = 16'hffff;
  rom[13121] = 16'hffff;
  rom[13122] = 16'hffff;
  rom[13123] = 16'hffff;
  rom[13124] = 16'hffff;
  rom[13125] = 16'hffff;
  rom[13126] = 16'hffff;
  rom[13127] = 16'hffff;
  rom[13128] = 16'hffff;
  rom[13129] = 16'hffff;
  rom[13130] = 16'hffff;
  rom[13131] = 16'hffff;
  rom[13132] = 16'hffff;
  rom[13133] = 16'hffff;
  rom[13134] = 16'hffff;
  rom[13135] = 16'hffff;
  rom[13136] = 16'hffff;
  rom[13137] = 16'hffff;
  rom[13138] = 16'hffde;
  rom[13139] = 16'h9c6e;
  rom[13140] = 16'hac2b;
  rom[13141] = 16'he56c;
  rom[13142] = 16'hfd6a;
  rom[13143] = 16'hfd48;
  rom[13144] = 16'hfd68;
  rom[13145] = 16'hfd48;
  rom[13146] = 16'hfd69;
  rom[13147] = 16'hfd68;
  rom[13148] = 16'hfd68;
  rom[13149] = 16'hfd47;
  rom[13150] = 16'hfd68;
  rom[13151] = 16'hf549;
  rom[13152] = 16'hf549;
  rom[13153] = 16'hed4a;
  rom[13154] = 16'h9306;
  rom[13155] = 16'hbd33;
  rom[13156] = 16'hffdf;
  rom[13157] = 16'hffff;
  rom[13158] = 16'hffff;
  rom[13159] = 16'hffff;
  rom[13160] = 16'hffff;
  rom[13161] = 16'hffff;
  rom[13162] = 16'hffff;
  rom[13163] = 16'hffff;
  rom[13164] = 16'hffff;
  rom[13165] = 16'hffff;
  rom[13166] = 16'hffff;
  rom[13167] = 16'hffff;
  rom[13168] = 16'hffff;
  rom[13169] = 16'hffff;
  rom[13170] = 16'hffff;
  rom[13171] = 16'hffff;
  rom[13172] = 16'hffff;
  rom[13173] = 16'hffff;
  rom[13174] = 16'hffff;
  rom[13175] = 16'hffff;
  rom[13176] = 16'hffff;
  rom[13177] = 16'hffff;
  rom[13178] = 16'hffff;
  rom[13179] = 16'hffff;
  rom[13180] = 16'hffff;
  rom[13181] = 16'hffff;
  rom[13182] = 16'hffff;
  rom[13183] = 16'hffff;
  rom[13184] = 16'hffff;
  rom[13185] = 16'hffff;
  rom[13186] = 16'hffff;
  rom[13187] = 16'hffff;
  rom[13188] = 16'hffff;
  rom[13189] = 16'hffff;
  rom[13190] = 16'hffff;
  rom[13191] = 16'hffff;
  rom[13192] = 16'hffff;
  rom[13193] = 16'hffff;
  rom[13194] = 16'hffff;
  rom[13195] = 16'hffff;
  rom[13196] = 16'hffff;
  rom[13197] = 16'hffff;
  rom[13198] = 16'hffff;
  rom[13199] = 16'hffff;
  rom[13200] = 16'hffff;
  rom[13201] = 16'hffff;
  rom[13202] = 16'hffff;
  rom[13203] = 16'hffff;
  rom[13204] = 16'hffff;
  rom[13205] = 16'hffff;
  rom[13206] = 16'hffff;
  rom[13207] = 16'hffff;
  rom[13208] = 16'hffff;
  rom[13209] = 16'hffff;
  rom[13210] = 16'hffff;
  rom[13211] = 16'hffff;
  rom[13212] = 16'hffff;
  rom[13213] = 16'hffff;
  rom[13214] = 16'hffff;
  rom[13215] = 16'hffff;
  rom[13216] = 16'hffff;
  rom[13217] = 16'hffff;
  rom[13218] = 16'hffff;
  rom[13219] = 16'hffff;
  rom[13220] = 16'hffff;
  rom[13221] = 16'hffff;
  rom[13222] = 16'hffff;
  rom[13223] = 16'hffff;
  rom[13224] = 16'hffff;
  rom[13225] = 16'hffff;
  rom[13226] = 16'hffff;
  rom[13227] = 16'hffff;
  rom[13228] = 16'hffff;
  rom[13229] = 16'hffff;
  rom[13230] = 16'hffff;
  rom[13231] = 16'hffff;
  rom[13232] = 16'hffff;
  rom[13233] = 16'hffff;
  rom[13234] = 16'hffff;
  rom[13235] = 16'hffff;
  rom[13236] = 16'hffff;
  rom[13237] = 16'hffff;
  rom[13238] = 16'hffff;
  rom[13239] = 16'hffff;
  rom[13240] = 16'hffdf;
  rom[13241] = 16'he698;
  rom[13242] = 16'h72c5;
  rom[13243] = 16'hdd2b;
  rom[13244] = 16'hf529;
  rom[13245] = 16'hf547;
  rom[13246] = 16'hf567;
  rom[13247] = 16'hf569;
  rom[13248] = 16'hf549;
  rom[13249] = 16'hfd68;
  rom[13250] = 16'hfd67;
  rom[13251] = 16'hfd69;
  rom[13252] = 16'he54b;
  rom[13253] = 16'hbccc;
  rom[13254] = 16'h8bab;
  rom[13255] = 16'hfffe;
  rom[13256] = 16'hffff;
  rom[13257] = 16'hffff;
  rom[13258] = 16'hffff;
  rom[13259] = 16'hffff;
  rom[13260] = 16'hffff;
  rom[13261] = 16'hffff;
  rom[13262] = 16'hffff;
  rom[13263] = 16'hffff;
  rom[13264] = 16'hffff;
  rom[13265] = 16'hffff;
  rom[13266] = 16'hffff;
  rom[13267] = 16'hffff;
  rom[13268] = 16'hffff;
  rom[13269] = 16'hffff;
  rom[13270] = 16'hffff;
  rom[13271] = 16'hffff;
  rom[13272] = 16'hffff;
  rom[13273] = 16'hffff;
  rom[13274] = 16'hffdf;
  rom[13275] = 16'hff9e;
  rom[13276] = 16'hdebb;
  rom[13277] = 16'hd659;
  rom[13278] = 16'hde9a;
  rom[13279] = 16'hf79e;
  rom[13280] = 16'hffff;
  rom[13281] = 16'hffff;
  rom[13282] = 16'hf7be;
  rom[13283] = 16'hffff;
  rom[13284] = 16'hffff;
  rom[13285] = 16'hffff;
  rom[13286] = 16'hffff;
  rom[13287] = 16'hffff;
  rom[13288] = 16'hffff;
  rom[13289] = 16'hffff;
  rom[13290] = 16'hffff;
  rom[13291] = 16'hffff;
  rom[13292] = 16'hffff;
  rom[13293] = 16'hffff;
  rom[13294] = 16'hffff;
  rom[13295] = 16'hffff;
  rom[13296] = 16'hffff;
  rom[13297] = 16'hffff;
  rom[13298] = 16'hffff;
  rom[13299] = 16'hffff;
  rom[13300] = 16'hffff;
  rom[13301] = 16'hffff;
  rom[13302] = 16'hffff;
  rom[13303] = 16'hffff;
  rom[13304] = 16'hffff;
  rom[13305] = 16'hffff;
  rom[13306] = 16'hffff;
  rom[13307] = 16'hffff;
  rom[13308] = 16'hffff;
  rom[13309] = 16'hffff;
  rom[13310] = 16'hffdf;
  rom[13311] = 16'hffff;
  rom[13312] = 16'hffbf;
  rom[13313] = 16'hffff;
  rom[13314] = 16'hffff;
  rom[13315] = 16'hef1c;
  rom[13316] = 16'hd679;
  rom[13317] = 16'hd699;
  rom[13318] = 16'hdedb;
  rom[13319] = 16'hffdf;
  rom[13320] = 16'hffff;
  rom[13321] = 16'hffff;
  rom[13322] = 16'hffdf;
  rom[13323] = 16'hffff;
  rom[13324] = 16'hffff;
  rom[13325] = 16'hffff;
  rom[13326] = 16'hffff;
  rom[13327] = 16'hffff;
  rom[13328] = 16'hffff;
  rom[13329] = 16'hffff;
  rom[13330] = 16'hffff;
  rom[13331] = 16'hffff;
  rom[13332] = 16'hffff;
  rom[13333] = 16'hffff;
  rom[13334] = 16'hffff;
  rom[13335] = 16'hffff;
  rom[13336] = 16'hffff;
  rom[13337] = 16'hffff;
  rom[13338] = 16'hffde;
  rom[13339] = 16'hce36;
  rom[13340] = 16'h8368;
  rom[13341] = 16'he54d;
  rom[13342] = 16'hed6a;
  rom[13343] = 16'hfd68;
  rom[13344] = 16'hfd47;
  rom[13345] = 16'hfd48;
  rom[13346] = 16'hf548;
  rom[13347] = 16'hfd68;
  rom[13348] = 16'hfd47;
  rom[13349] = 16'hfd68;
  rom[13350] = 16'hf547;
  rom[13351] = 16'hf549;
  rom[13352] = 16'hfd29;
  rom[13353] = 16'hf54b;
  rom[13354] = 16'h9305;
  rom[13355] = 16'hbcf3;
  rom[13356] = 16'hffbf;
  rom[13357] = 16'hffff;
  rom[13358] = 16'hffff;
  rom[13359] = 16'hffff;
  rom[13360] = 16'hffff;
  rom[13361] = 16'hffff;
  rom[13362] = 16'hffff;
  rom[13363] = 16'hffff;
  rom[13364] = 16'hffff;
  rom[13365] = 16'hffff;
  rom[13366] = 16'hffff;
  rom[13367] = 16'hffff;
  rom[13368] = 16'hffff;
  rom[13369] = 16'hffff;
  rom[13370] = 16'hffff;
  rom[13371] = 16'hffff;
  rom[13372] = 16'hffff;
  rom[13373] = 16'hffff;
  rom[13374] = 16'hffff;
  rom[13375] = 16'hffff;
  rom[13376] = 16'hffff;
  rom[13377] = 16'hffff;
  rom[13378] = 16'hffff;
  rom[13379] = 16'hffff;
  rom[13380] = 16'hffff;
  rom[13381] = 16'hffff;
  rom[13382] = 16'hffff;
  rom[13383] = 16'hffff;
  rom[13384] = 16'hffff;
  rom[13385] = 16'hffff;
  rom[13386] = 16'hffff;
  rom[13387] = 16'hffff;
  rom[13388] = 16'hffff;
  rom[13389] = 16'hffff;
  rom[13390] = 16'hffff;
  rom[13391] = 16'hffff;
  rom[13392] = 16'hffff;
  rom[13393] = 16'hffff;
  rom[13394] = 16'hffff;
  rom[13395] = 16'hffff;
  rom[13396] = 16'hffff;
  rom[13397] = 16'hffff;
  rom[13398] = 16'hffff;
  rom[13399] = 16'hffff;
  rom[13400] = 16'hffff;
  rom[13401] = 16'hffff;
  rom[13402] = 16'hffff;
  rom[13403] = 16'hffff;
  rom[13404] = 16'hffff;
  rom[13405] = 16'hffff;
  rom[13406] = 16'hffff;
  rom[13407] = 16'hffff;
  rom[13408] = 16'hffff;
  rom[13409] = 16'hffff;
  rom[13410] = 16'hffff;
  rom[13411] = 16'hffff;
  rom[13412] = 16'hffff;
  rom[13413] = 16'hffff;
  rom[13414] = 16'hffff;
  rom[13415] = 16'hffff;
  rom[13416] = 16'hffff;
  rom[13417] = 16'hffff;
  rom[13418] = 16'hffff;
  rom[13419] = 16'hffff;
  rom[13420] = 16'hffff;
  rom[13421] = 16'hffff;
  rom[13422] = 16'hffff;
  rom[13423] = 16'hffff;
  rom[13424] = 16'hffff;
  rom[13425] = 16'hffff;
  rom[13426] = 16'hffff;
  rom[13427] = 16'hffff;
  rom[13428] = 16'hffff;
  rom[13429] = 16'hffff;
  rom[13430] = 16'hffff;
  rom[13431] = 16'hffff;
  rom[13432] = 16'hffff;
  rom[13433] = 16'hffff;
  rom[13434] = 16'hffff;
  rom[13435] = 16'hffff;
  rom[13436] = 16'hffff;
  rom[13437] = 16'hffff;
  rom[13438] = 16'hffff;
  rom[13439] = 16'hffdf;
  rom[13440] = 16'hffff;
  rom[13441] = 16'hcdb5;
  rom[13442] = 16'h93a9;
  rom[13443] = 16'hdd6c;
  rom[13444] = 16'hfdaa;
  rom[13445] = 16'hf527;
  rom[13446] = 16'hfd88;
  rom[13447] = 16'hf548;
  rom[13448] = 16'hfd6a;
  rom[13449] = 16'hfd49;
  rom[13450] = 16'hfd69;
  rom[13451] = 16'hfd49;
  rom[13452] = 16'he5ad;
  rom[13453] = 16'h9387;
  rom[13454] = 16'hc593;
  rom[13455] = 16'hffde;
  rom[13456] = 16'hffff;
  rom[13457] = 16'hffff;
  rom[13458] = 16'hffff;
  rom[13459] = 16'hffff;
  rom[13460] = 16'hffff;
  rom[13461] = 16'hffff;
  rom[13462] = 16'hffff;
  rom[13463] = 16'hffff;
  rom[13464] = 16'hffff;
  rom[13465] = 16'hffff;
  rom[13466] = 16'hffff;
  rom[13467] = 16'hffff;
  rom[13468] = 16'hffff;
  rom[13469] = 16'hffff;
  rom[13470] = 16'hffff;
  rom[13471] = 16'hffff;
  rom[13472] = 16'hffdf;
  rom[13473] = 16'hce18;
  rom[13474] = 16'h7bae;
  rom[13475] = 16'h41e8;
  rom[13476] = 16'h3166;
  rom[13477] = 16'h2945;
  rom[13478] = 16'h39a6;
  rom[13479] = 16'h4248;
  rom[13480] = 16'h6b2d;
  rom[13481] = 16'hc5f8;
  rom[13482] = 16'hf77e;
  rom[13483] = 16'hffdf;
  rom[13484] = 16'hffff;
  rom[13485] = 16'hffff;
  rom[13486] = 16'hffff;
  rom[13487] = 16'hffff;
  rom[13488] = 16'hffff;
  rom[13489] = 16'hffff;
  rom[13490] = 16'hffff;
  rom[13491] = 16'hffff;
  rom[13492] = 16'hffff;
  rom[13493] = 16'hffff;
  rom[13494] = 16'hffff;
  rom[13495] = 16'hffff;
  rom[13496] = 16'hffff;
  rom[13497] = 16'hffff;
  rom[13498] = 16'hffff;
  rom[13499] = 16'hffff;
  rom[13500] = 16'hffff;
  rom[13501] = 16'hffff;
  rom[13502] = 16'hffff;
  rom[13503] = 16'hffff;
  rom[13504] = 16'hffff;
  rom[13505] = 16'hffff;
  rom[13506] = 16'hffff;
  rom[13507] = 16'hffff;
  rom[13508] = 16'hffff;
  rom[13509] = 16'hffff;
  rom[13510] = 16'hffff;
  rom[13511] = 16'hffbf;
  rom[13512] = 16'hef3d;
  rom[13513] = 16'h9492;
  rom[13514] = 16'h5aaa;
  rom[13515] = 16'h39c6;
  rom[13516] = 16'h3165;
  rom[13517] = 16'h2124;
  rom[13518] = 16'h39a6;
  rom[13519] = 16'h5aaa;
  rom[13520] = 16'h9cd3;
  rom[13521] = 16'hf7be;
  rom[13522] = 16'hffff;
  rom[13523] = 16'hffff;
  rom[13524] = 16'hffff;
  rom[13525] = 16'hffff;
  rom[13526] = 16'hffff;
  rom[13527] = 16'hffff;
  rom[13528] = 16'hffff;
  rom[13529] = 16'hffff;
  rom[13530] = 16'hffff;
  rom[13531] = 16'hffff;
  rom[13532] = 16'hffff;
  rom[13533] = 16'hffff;
  rom[13534] = 16'hffff;
  rom[13535] = 16'hffff;
  rom[13536] = 16'hffff;
  rom[13537] = 16'hffff;
  rom[13538] = 16'hffff;
  rom[13539] = 16'hef3b;
  rom[13540] = 16'h8baa;
  rom[13541] = 16'hbc6a;
  rom[13542] = 16'hf5ab;
  rom[13543] = 16'hfd68;
  rom[13544] = 16'hfd48;
  rom[13545] = 16'hfd69;
  rom[13546] = 16'hfd68;
  rom[13547] = 16'hfd48;
  rom[13548] = 16'hfd69;
  rom[13549] = 16'hf528;
  rom[13550] = 16'hfd69;
  rom[13551] = 16'hf549;
  rom[13552] = 16'hfd4a;
  rom[13553] = 16'hf52b;
  rom[13554] = 16'h9b26;
  rom[13555] = 16'hb4f3;
  rom[13556] = 16'hffdf;
  rom[13557] = 16'hffff;
  rom[13558] = 16'hffff;
  rom[13559] = 16'hffff;
  rom[13560] = 16'hffff;
  rom[13561] = 16'hffff;
  rom[13562] = 16'hffff;
  rom[13563] = 16'hffff;
  rom[13564] = 16'hffff;
  rom[13565] = 16'hffff;
  rom[13566] = 16'hffff;
  rom[13567] = 16'hffff;
  rom[13568] = 16'hffff;
  rom[13569] = 16'hffff;
  rom[13570] = 16'hffff;
  rom[13571] = 16'hffff;
  rom[13572] = 16'hffff;
  rom[13573] = 16'hffff;
  rom[13574] = 16'hffff;
  rom[13575] = 16'hffff;
  rom[13576] = 16'hffff;
  rom[13577] = 16'hffff;
  rom[13578] = 16'hffff;
  rom[13579] = 16'hffff;
  rom[13580] = 16'hffff;
  rom[13581] = 16'hffff;
  rom[13582] = 16'hffff;
  rom[13583] = 16'hffff;
  rom[13584] = 16'hffff;
  rom[13585] = 16'hffff;
  rom[13586] = 16'hffff;
  rom[13587] = 16'hffff;
  rom[13588] = 16'hffff;
  rom[13589] = 16'hffff;
  rom[13590] = 16'hffff;
  rom[13591] = 16'hffff;
  rom[13592] = 16'hffff;
  rom[13593] = 16'hffff;
  rom[13594] = 16'hffff;
  rom[13595] = 16'hffff;
  rom[13596] = 16'hffff;
  rom[13597] = 16'hffff;
  rom[13598] = 16'hffff;
  rom[13599] = 16'hffff;
  rom[13600] = 16'hffff;
  rom[13601] = 16'hffff;
  rom[13602] = 16'hffff;
  rom[13603] = 16'hffff;
  rom[13604] = 16'hffff;
  rom[13605] = 16'hffff;
  rom[13606] = 16'hffff;
  rom[13607] = 16'hffff;
  rom[13608] = 16'hffff;
  rom[13609] = 16'hffff;
  rom[13610] = 16'hffff;
  rom[13611] = 16'hffff;
  rom[13612] = 16'hffff;
  rom[13613] = 16'hffff;
  rom[13614] = 16'hffff;
  rom[13615] = 16'hffff;
  rom[13616] = 16'hffff;
  rom[13617] = 16'hffff;
  rom[13618] = 16'hffff;
  rom[13619] = 16'hffff;
  rom[13620] = 16'hffff;
  rom[13621] = 16'hffff;
  rom[13622] = 16'hffff;
  rom[13623] = 16'hffff;
  rom[13624] = 16'hffff;
  rom[13625] = 16'hffff;
  rom[13626] = 16'hffff;
  rom[13627] = 16'hffff;
  rom[13628] = 16'hffff;
  rom[13629] = 16'hffff;
  rom[13630] = 16'hffff;
  rom[13631] = 16'hffff;
  rom[13632] = 16'hffff;
  rom[13633] = 16'hffff;
  rom[13634] = 16'hffff;
  rom[13635] = 16'hffff;
  rom[13636] = 16'hfffe;
  rom[13637] = 16'hffff;
  rom[13638] = 16'hffdf;
  rom[13639] = 16'hffff;
  rom[13640] = 16'hffdf;
  rom[13641] = 16'ha44e;
  rom[13642] = 16'hac09;
  rom[13643] = 16'hed4b;
  rom[13644] = 16'hed27;
  rom[13645] = 16'hf548;
  rom[13646] = 16'hfd48;
  rom[13647] = 16'hfd48;
  rom[13648] = 16'hfd28;
  rom[13649] = 16'hfd49;
  rom[13650] = 16'hfd48;
  rom[13651] = 16'hfd89;
  rom[13652] = 16'hcd4b;
  rom[13653] = 16'h7b27;
  rom[13654] = 16'he6d8;
  rom[13655] = 16'hffdf;
  rom[13656] = 16'hfffe;
  rom[13657] = 16'hffff;
  rom[13658] = 16'hffff;
  rom[13659] = 16'hffff;
  rom[13660] = 16'hffff;
  rom[13661] = 16'hffff;
  rom[13662] = 16'hffff;
  rom[13663] = 16'hffff;
  rom[13664] = 16'hffff;
  rom[13665] = 16'hffff;
  rom[13666] = 16'hffff;
  rom[13667] = 16'hffff;
  rom[13668] = 16'hffff;
  rom[13669] = 16'hffdf;
  rom[13670] = 16'hffff;
  rom[13671] = 16'hffff;
  rom[13672] = 16'hf77d;
  rom[13673] = 16'h83f0;
  rom[13674] = 16'h2924;
  rom[13675] = 16'h5aab;
  rom[13676] = 16'h83f0;
  rom[13677] = 16'h9492;
  rom[13678] = 16'h83f0;
  rom[13679] = 16'h5289;
  rom[13680] = 16'h2144;
  rom[13681] = 16'h2924;
  rom[13682] = 16'h4a48;
  rom[13683] = 16'h9cb2;
  rom[13684] = 16'he71c;
  rom[13685] = 16'hffff;
  rom[13686] = 16'hffff;
  rom[13687] = 16'hffff;
  rom[13688] = 16'hffff;
  rom[13689] = 16'hffff;
  rom[13690] = 16'hffff;
  rom[13691] = 16'hffff;
  rom[13692] = 16'hffff;
  rom[13693] = 16'hffff;
  rom[13694] = 16'hffff;
  rom[13695] = 16'hffff;
  rom[13696] = 16'hffff;
  rom[13697] = 16'hffff;
  rom[13698] = 16'hffff;
  rom[13699] = 16'hffff;
  rom[13700] = 16'hffff;
  rom[13701] = 16'hffff;
  rom[13702] = 16'hffff;
  rom[13703] = 16'hffff;
  rom[13704] = 16'hffff;
  rom[13705] = 16'hffff;
  rom[13706] = 16'hffff;
  rom[13707] = 16'hffff;
  rom[13708] = 16'hffff;
  rom[13709] = 16'hffdf;
  rom[13710] = 16'hbdf7;
  rom[13711] = 16'h734d;
  rom[13712] = 16'h2965;
  rom[13713] = 16'h2104;
  rom[13714] = 16'h39c6;
  rom[13715] = 16'h6b4d;
  rom[13716] = 16'h8c51;
  rom[13717] = 16'h9492;
  rom[13718] = 16'h738e;
  rom[13719] = 16'h49e7;
  rom[13720] = 16'h39a6;
  rom[13721] = 16'hd6ba;
  rom[13722] = 16'hffdf;
  rom[13723] = 16'hffff;
  rom[13724] = 16'hffdf;
  rom[13725] = 16'hffff;
  rom[13726] = 16'hffff;
  rom[13727] = 16'hffff;
  rom[13728] = 16'hffff;
  rom[13729] = 16'hffff;
  rom[13730] = 16'hffff;
  rom[13731] = 16'hffff;
  rom[13732] = 16'hffff;
  rom[13733] = 16'hffff;
  rom[13734] = 16'hffff;
  rom[13735] = 16'hffff;
  rom[13736] = 16'hffff;
  rom[13737] = 16'hffff;
  rom[13738] = 16'hffff;
  rom[13739] = 16'hffde;
  rom[13740] = 16'h946e;
  rom[13741] = 16'h93a9;
  rom[13742] = 16'he56b;
  rom[13743] = 16'hf588;
  rom[13744] = 16'hfd48;
  rom[13745] = 16'hfd49;
  rom[13746] = 16'hfd08;
  rom[13747] = 16'hfd48;
  rom[13748] = 16'hf529;
  rom[13749] = 16'hf569;
  rom[13750] = 16'hf548;
  rom[13751] = 16'hfd48;
  rom[13752] = 16'hf528;
  rom[13753] = 16'hed4b;
  rom[13754] = 16'h8ae6;
  rom[13755] = 16'hbd33;
  rom[13756] = 16'hffde;
  rom[13757] = 16'hffff;
  rom[13758] = 16'hffff;
  rom[13759] = 16'hffff;
  rom[13760] = 16'hffff;
  rom[13761] = 16'hffff;
  rom[13762] = 16'hffff;
  rom[13763] = 16'hffff;
  rom[13764] = 16'hffff;
  rom[13765] = 16'hffff;
  rom[13766] = 16'hffff;
  rom[13767] = 16'hffff;
  rom[13768] = 16'hffff;
  rom[13769] = 16'hffff;
  rom[13770] = 16'hffff;
  rom[13771] = 16'hffff;
  rom[13772] = 16'hffff;
  rom[13773] = 16'hffff;
  rom[13774] = 16'hffff;
  rom[13775] = 16'hffff;
  rom[13776] = 16'hffff;
  rom[13777] = 16'hffff;
  rom[13778] = 16'hffff;
  rom[13779] = 16'hffff;
  rom[13780] = 16'hffff;
  rom[13781] = 16'hffff;
  rom[13782] = 16'hffff;
  rom[13783] = 16'hffff;
  rom[13784] = 16'hffff;
  rom[13785] = 16'hffff;
  rom[13786] = 16'hffff;
  rom[13787] = 16'hffff;
  rom[13788] = 16'hffff;
  rom[13789] = 16'hffff;
  rom[13790] = 16'hffff;
  rom[13791] = 16'hffff;
  rom[13792] = 16'hffff;
  rom[13793] = 16'hffff;
  rom[13794] = 16'hffff;
  rom[13795] = 16'hffff;
  rom[13796] = 16'hffff;
  rom[13797] = 16'hffff;
  rom[13798] = 16'hffff;
  rom[13799] = 16'hffff;
  rom[13800] = 16'hffff;
  rom[13801] = 16'hffff;
  rom[13802] = 16'hffff;
  rom[13803] = 16'hffff;
  rom[13804] = 16'hffff;
  rom[13805] = 16'hffff;
  rom[13806] = 16'hffff;
  rom[13807] = 16'hffff;
  rom[13808] = 16'hffff;
  rom[13809] = 16'hffff;
  rom[13810] = 16'hffff;
  rom[13811] = 16'hffff;
  rom[13812] = 16'hffff;
  rom[13813] = 16'hffff;
  rom[13814] = 16'hffff;
  rom[13815] = 16'hffff;
  rom[13816] = 16'hffff;
  rom[13817] = 16'hffff;
  rom[13818] = 16'hffff;
  rom[13819] = 16'hffff;
  rom[13820] = 16'hffff;
  rom[13821] = 16'hffff;
  rom[13822] = 16'hffff;
  rom[13823] = 16'hffff;
  rom[13824] = 16'hffff;
  rom[13825] = 16'hffff;
  rom[13826] = 16'hffff;
  rom[13827] = 16'hffff;
  rom[13828] = 16'hffff;
  rom[13829] = 16'hffff;
  rom[13830] = 16'hffff;
  rom[13831] = 16'hffff;
  rom[13832] = 16'hffff;
  rom[13833] = 16'hffff;
  rom[13834] = 16'hffff;
  rom[13835] = 16'hffff;
  rom[13836] = 16'hffdf;
  rom[13837] = 16'hffff;
  rom[13838] = 16'hffff;
  rom[13839] = 16'hffff;
  rom[13840] = 16'hef3c;
  rom[13841] = 16'h93ab;
  rom[13842] = 16'hc4ab;
  rom[13843] = 16'hfdec;
  rom[13844] = 16'hfd68;
  rom[13845] = 16'hfd68;
  rom[13846] = 16'hf528;
  rom[13847] = 16'hfd28;
  rom[13848] = 16'hfd6a;
  rom[13849] = 16'hfd28;
  rom[13850] = 16'hfd89;
  rom[13851] = 16'hed48;
  rom[13852] = 16'hc4eb;
  rom[13853] = 16'h7328;
  rom[13854] = 16'hf73c;
  rom[13855] = 16'hffff;
  rom[13856] = 16'hffff;
  rom[13857] = 16'hffff;
  rom[13858] = 16'hffff;
  rom[13859] = 16'hffff;
  rom[13860] = 16'hffff;
  rom[13861] = 16'hffff;
  rom[13862] = 16'hffff;
  rom[13863] = 16'hffff;
  rom[13864] = 16'hffff;
  rom[13865] = 16'hffff;
  rom[13866] = 16'hffff;
  rom[13867] = 16'hffff;
  rom[13868] = 16'hffff;
  rom[13869] = 16'hffff;
  rom[13870] = 16'hffff;
  rom[13871] = 16'hffbf;
  rom[13872] = 16'hffff;
  rom[13873] = 16'hef5d;
  rom[13874] = 16'hffff;
  rom[13875] = 16'hffbf;
  rom[13876] = 16'hffff;
  rom[13877] = 16'hffff;
  rom[13878] = 16'hffff;
  rom[13879] = 16'hf79e;
  rom[13880] = 16'hef5d;
  rom[13881] = 16'h7bcf;
  rom[13882] = 16'h3166;
  rom[13883] = 16'h18c2;
  rom[13884] = 16'h4208;
  rom[13885] = 16'hb596;
  rom[13886] = 16'hffff;
  rom[13887] = 16'hffff;
  rom[13888] = 16'hffff;
  rom[13889] = 16'hffff;
  rom[13890] = 16'hffff;
  rom[13891] = 16'hffff;
  rom[13892] = 16'hffff;
  rom[13893] = 16'hffff;
  rom[13894] = 16'hffff;
  rom[13895] = 16'hffff;
  rom[13896] = 16'hffff;
  rom[13897] = 16'hffff;
  rom[13898] = 16'hffff;
  rom[13899] = 16'hffff;
  rom[13900] = 16'hffff;
  rom[13901] = 16'hffff;
  rom[13902] = 16'hffff;
  rom[13903] = 16'hffff;
  rom[13904] = 16'hffff;
  rom[13905] = 16'hffff;
  rom[13906] = 16'hffff;
  rom[13907] = 16'hffff;
  rom[13908] = 16'hf77d;
  rom[13909] = 16'h73ce;
  rom[13910] = 16'h18a2;
  rom[13911] = 16'h2124;
  rom[13912] = 16'h5a8a;
  rom[13913] = 16'hc638;
  rom[13914] = 16'hff9e;
  rom[13915] = 16'hffff;
  rom[13916] = 16'hffff;
  rom[13917] = 16'hffff;
  rom[13918] = 16'hffff;
  rom[13919] = 16'hffbe;
  rom[13920] = 16'hffdf;
  rom[13921] = 16'hffff;
  rom[13922] = 16'hffff;
  rom[13923] = 16'hffff;
  rom[13924] = 16'hffdf;
  rom[13925] = 16'hffff;
  rom[13926] = 16'hffff;
  rom[13927] = 16'hffff;
  rom[13928] = 16'hffff;
  rom[13929] = 16'hffff;
  rom[13930] = 16'hffff;
  rom[13931] = 16'hffff;
  rom[13932] = 16'hffff;
  rom[13933] = 16'hffff;
  rom[13934] = 16'hffff;
  rom[13935] = 16'hffff;
  rom[13936] = 16'hffff;
  rom[13937] = 16'hffff;
  rom[13938] = 16'hffff;
  rom[13939] = 16'hffff;
  rom[13940] = 16'hcdf5;
  rom[13941] = 16'h9c0b;
  rom[13942] = 16'he56c;
  rom[13943] = 16'hf547;
  rom[13944] = 16'hfd49;
  rom[13945] = 16'hfd49;
  rom[13946] = 16'hfd89;
  rom[13947] = 16'hfd28;
  rom[13948] = 16'hfd4a;
  rom[13949] = 16'hf569;
  rom[13950] = 16'hfd69;
  rom[13951] = 16'hfd28;
  rom[13952] = 16'hfd49;
  rom[13953] = 16'he52b;
  rom[13954] = 16'h8ae6;
  rom[13955] = 16'hbd75;
  rom[13956] = 16'hffff;
  rom[13957] = 16'hffff;
  rom[13958] = 16'hffff;
  rom[13959] = 16'hffff;
  rom[13960] = 16'hffff;
  rom[13961] = 16'hffff;
  rom[13962] = 16'hffff;
  rom[13963] = 16'hffff;
  rom[13964] = 16'hffff;
  rom[13965] = 16'hffff;
  rom[13966] = 16'hffff;
  rom[13967] = 16'hffff;
  rom[13968] = 16'hffff;
  rom[13969] = 16'hffff;
  rom[13970] = 16'hffff;
  rom[13971] = 16'hffff;
  rom[13972] = 16'hffff;
  rom[13973] = 16'hffff;
  rom[13974] = 16'hffff;
  rom[13975] = 16'hffff;
  rom[13976] = 16'hffff;
  rom[13977] = 16'hffff;
  rom[13978] = 16'hffff;
  rom[13979] = 16'hffff;
  rom[13980] = 16'hffff;
  rom[13981] = 16'hffff;
  rom[13982] = 16'hffff;
  rom[13983] = 16'hffff;
  rom[13984] = 16'hffff;
  rom[13985] = 16'hffff;
  rom[13986] = 16'hffff;
  rom[13987] = 16'hffff;
  rom[13988] = 16'hffff;
  rom[13989] = 16'hffff;
  rom[13990] = 16'hffff;
  rom[13991] = 16'hffff;
  rom[13992] = 16'hffff;
  rom[13993] = 16'hffff;
  rom[13994] = 16'hffff;
  rom[13995] = 16'hffff;
  rom[13996] = 16'hffff;
  rom[13997] = 16'hffff;
  rom[13998] = 16'hffff;
  rom[13999] = 16'hffff;
  rom[14000] = 16'hffff;
  rom[14001] = 16'hffff;
  rom[14002] = 16'hffff;
  rom[14003] = 16'hffff;
  rom[14004] = 16'hffff;
  rom[14005] = 16'hffff;
  rom[14006] = 16'hffff;
  rom[14007] = 16'hffff;
  rom[14008] = 16'hffff;
  rom[14009] = 16'hffff;
  rom[14010] = 16'hffff;
  rom[14011] = 16'hffff;
  rom[14012] = 16'hffff;
  rom[14013] = 16'hffff;
  rom[14014] = 16'hffff;
  rom[14015] = 16'hffff;
  rom[14016] = 16'hffff;
  rom[14017] = 16'hffff;
  rom[14018] = 16'hffff;
  rom[14019] = 16'hffff;
  rom[14020] = 16'hffff;
  rom[14021] = 16'hffff;
  rom[14022] = 16'hffff;
  rom[14023] = 16'hffff;
  rom[14024] = 16'hffff;
  rom[14025] = 16'hffff;
  rom[14026] = 16'hffff;
  rom[14027] = 16'hffff;
  rom[14028] = 16'hffff;
  rom[14029] = 16'hffff;
  rom[14030] = 16'hffff;
  rom[14031] = 16'hffff;
  rom[14032] = 16'hffff;
  rom[14033] = 16'hffff;
  rom[14034] = 16'hffff;
  rom[14035] = 16'hffff;
  rom[14036] = 16'hffdf;
  rom[14037] = 16'hffff;
  rom[14038] = 16'hf7df;
  rom[14039] = 16'hffff;
  rom[14040] = 16'hde99;
  rom[14041] = 16'h6a24;
  rom[14042] = 16'hdd2c;
  rom[14043] = 16'hed08;
  rom[14044] = 16'hfd48;
  rom[14045] = 16'hfd68;
  rom[14046] = 16'hfd88;
  rom[14047] = 16'hfd69;
  rom[14048] = 16'hfd28;
  rom[14049] = 16'hfd69;
  rom[14050] = 16'hed47;
  rom[14051] = 16'hed89;
  rom[14052] = 16'ha409;
  rom[14053] = 16'h942f;
  rom[14054] = 16'hffbe;
  rom[14055] = 16'hffff;
  rom[14056] = 16'hffff;
  rom[14057] = 16'hffff;
  rom[14058] = 16'hffff;
  rom[14059] = 16'hffff;
  rom[14060] = 16'hffff;
  rom[14061] = 16'hffff;
  rom[14062] = 16'hffff;
  rom[14063] = 16'hffff;
  rom[14064] = 16'hffff;
  rom[14065] = 16'hffff;
  rom[14066] = 16'hffff;
  rom[14067] = 16'hffff;
  rom[14068] = 16'hffff;
  rom[14069] = 16'hffff;
  rom[14070] = 16'hffff;
  rom[14071] = 16'hffff;
  rom[14072] = 16'hffff;
  rom[14073] = 16'hffff;
  rom[14074] = 16'hffdf;
  rom[14075] = 16'hffff;
  rom[14076] = 16'hffdf;
  rom[14077] = 16'hffff;
  rom[14078] = 16'hffdf;
  rom[14079] = 16'hffff;
  rom[14080] = 16'hffdf;
  rom[14081] = 16'hffff;
  rom[14082] = 16'he6fb;
  rom[14083] = 16'h8c71;
  rom[14084] = 16'h31a6;
  rom[14085] = 16'h2965;
  rom[14086] = 16'h8410;
  rom[14087] = 16'hef3c;
  rom[14088] = 16'hffdf;
  rom[14089] = 16'hffff;
  rom[14090] = 16'hffff;
  rom[14091] = 16'hffff;
  rom[14092] = 16'hffff;
  rom[14093] = 16'hffff;
  rom[14094] = 16'hffff;
  rom[14095] = 16'hffff;
  rom[14096] = 16'hffff;
  rom[14097] = 16'hffff;
  rom[14098] = 16'hffff;
  rom[14099] = 16'hffff;
  rom[14100] = 16'hffff;
  rom[14101] = 16'hffff;
  rom[14102] = 16'hffff;
  rom[14103] = 16'hffff;
  rom[14104] = 16'hffde;
  rom[14105] = 16'hffff;
  rom[14106] = 16'hf77d;
  rom[14107] = 16'hbdd6;
  rom[14108] = 16'h4a28;
  rom[14109] = 16'h2944;
  rom[14110] = 16'h52a9;
  rom[14111] = 16'hbdb6;
  rom[14112] = 16'hffff;
  rom[14113] = 16'hffdf;
  rom[14114] = 16'hffdf;
  rom[14115] = 16'hffff;
  rom[14116] = 16'hffff;
  rom[14117] = 16'hffff;
  rom[14118] = 16'hffff;
  rom[14119] = 16'hffff;
  rom[14120] = 16'hffdf;
  rom[14121] = 16'hffff;
  rom[14122] = 16'hffff;
  rom[14123] = 16'hffff;
  rom[14124] = 16'hffff;
  rom[14125] = 16'hffff;
  rom[14126] = 16'hffff;
  rom[14127] = 16'hffff;
  rom[14128] = 16'hffff;
  rom[14129] = 16'hffff;
  rom[14130] = 16'hffff;
  rom[14131] = 16'hffff;
  rom[14132] = 16'hffff;
  rom[14133] = 16'hffff;
  rom[14134] = 16'hffff;
  rom[14135] = 16'hffff;
  rom[14136] = 16'hffff;
  rom[14137] = 16'hffff;
  rom[14138] = 16'hffff;
  rom[14139] = 16'hffff;
  rom[14140] = 16'he6fa;
  rom[14141] = 16'h72c7;
  rom[14142] = 16'hc4ca;
  rom[14143] = 16'hfda9;
  rom[14144] = 16'hfd48;
  rom[14145] = 16'hf528;
  rom[14146] = 16'hfd48;
  rom[14147] = 16'hfd48;
  rom[14148] = 16'hfd29;
  rom[14149] = 16'hfd49;
  rom[14150] = 16'hf548;
  rom[14151] = 16'hfd27;
  rom[14152] = 16'hf549;
  rom[14153] = 16'hdd2b;
  rom[14154] = 16'h7ac5;
  rom[14155] = 16'hde38;
  rom[14156] = 16'hffdf;
  rom[14157] = 16'hffff;
  rom[14158] = 16'hffff;
  rom[14159] = 16'hffff;
  rom[14160] = 16'hffff;
  rom[14161] = 16'hffff;
  rom[14162] = 16'hffff;
  rom[14163] = 16'hffff;
  rom[14164] = 16'hffff;
  rom[14165] = 16'hffff;
  rom[14166] = 16'hffff;
  rom[14167] = 16'hffff;
  rom[14168] = 16'hffff;
  rom[14169] = 16'hffff;
  rom[14170] = 16'hffff;
  rom[14171] = 16'hffff;
  rom[14172] = 16'hffff;
  rom[14173] = 16'hffff;
  rom[14174] = 16'hffff;
  rom[14175] = 16'hffff;
  rom[14176] = 16'hffff;
  rom[14177] = 16'hffff;
  rom[14178] = 16'hffff;
  rom[14179] = 16'hffff;
  rom[14180] = 16'hffff;
  rom[14181] = 16'hffff;
  rom[14182] = 16'hffff;
  rom[14183] = 16'hffff;
  rom[14184] = 16'hffff;
  rom[14185] = 16'hffff;
  rom[14186] = 16'hffff;
  rom[14187] = 16'hffff;
  rom[14188] = 16'hffff;
  rom[14189] = 16'hffff;
  rom[14190] = 16'hffff;
  rom[14191] = 16'hffff;
  rom[14192] = 16'hffff;
  rom[14193] = 16'hffff;
  rom[14194] = 16'hffff;
  rom[14195] = 16'hffff;
  rom[14196] = 16'hffff;
  rom[14197] = 16'hffff;
  rom[14198] = 16'hffff;
  rom[14199] = 16'hffff;
  rom[14200] = 16'hffff;
  rom[14201] = 16'hffff;
  rom[14202] = 16'hffff;
  rom[14203] = 16'hffff;
  rom[14204] = 16'hffff;
  rom[14205] = 16'hffff;
  rom[14206] = 16'hffff;
  rom[14207] = 16'hffff;
  rom[14208] = 16'hffff;
  rom[14209] = 16'hffff;
  rom[14210] = 16'hffff;
  rom[14211] = 16'hffff;
  rom[14212] = 16'hffff;
  rom[14213] = 16'hffff;
  rom[14214] = 16'hffff;
  rom[14215] = 16'hffff;
  rom[14216] = 16'hffff;
  rom[14217] = 16'hffff;
  rom[14218] = 16'hffff;
  rom[14219] = 16'hffff;
  rom[14220] = 16'hffff;
  rom[14221] = 16'hffff;
  rom[14222] = 16'hffff;
  rom[14223] = 16'hffff;
  rom[14224] = 16'hffff;
  rom[14225] = 16'hffff;
  rom[14226] = 16'hffff;
  rom[14227] = 16'hffff;
  rom[14228] = 16'hffff;
  rom[14229] = 16'hffff;
  rom[14230] = 16'hffff;
  rom[14231] = 16'hffff;
  rom[14232] = 16'hffff;
  rom[14233] = 16'hffff;
  rom[14234] = 16'hffff;
  rom[14235] = 16'hffff;
  rom[14236] = 16'hffff;
  rom[14237] = 16'hffff;
  rom[14238] = 16'hffff;
  rom[14239] = 16'hffff;
  rom[14240] = 16'hb532;
  rom[14241] = 16'h7ac5;
  rom[14242] = 16'he54c;
  rom[14243] = 16'hfd29;
  rom[14244] = 16'hfd49;
  rom[14245] = 16'hed06;
  rom[14246] = 16'hf548;
  rom[14247] = 16'hfd48;
  rom[14248] = 16'hfd49;
  rom[14249] = 16'hfd68;
  rom[14250] = 16'hfda8;
  rom[14251] = 16'hed89;
  rom[14252] = 16'h9389;
  rom[14253] = 16'hbd75;
  rom[14254] = 16'hffdf;
  rom[14255] = 16'hffff;
  rom[14256] = 16'hffff;
  rom[14257] = 16'hffff;
  rom[14258] = 16'hffff;
  rom[14259] = 16'hffff;
  rom[14260] = 16'hffff;
  rom[14261] = 16'hffff;
  rom[14262] = 16'hffff;
  rom[14263] = 16'hffff;
  rom[14264] = 16'hffff;
  rom[14265] = 16'hffff;
  rom[14266] = 16'hffff;
  rom[14267] = 16'hffff;
  rom[14268] = 16'hffff;
  rom[14269] = 16'hffff;
  rom[14270] = 16'hffff;
  rom[14271] = 16'hffff;
  rom[14272] = 16'hffff;
  rom[14273] = 16'hffff;
  rom[14274] = 16'hffff;
  rom[14275] = 16'hffff;
  rom[14276] = 16'hffff;
  rom[14277] = 16'hffff;
  rom[14278] = 16'hffff;
  rom[14279] = 16'hffdf;
  rom[14280] = 16'hffff;
  rom[14281] = 16'hffff;
  rom[14282] = 16'hffff;
  rom[14283] = 16'hffdf;
  rom[14284] = 16'hce59;
  rom[14285] = 16'h5aeb;
  rom[14286] = 16'h18c3;
  rom[14287] = 16'h6b4d;
  rom[14288] = 16'hf77e;
  rom[14289] = 16'hffff;
  rom[14290] = 16'hffff;
  rom[14291] = 16'hffff;
  rom[14292] = 16'hffff;
  rom[14293] = 16'hffff;
  rom[14294] = 16'hffff;
  rom[14295] = 16'hffff;
  rom[14296] = 16'hffff;
  rom[14297] = 16'hffff;
  rom[14298] = 16'hffff;
  rom[14299] = 16'hffff;
  rom[14300] = 16'hffff;
  rom[14301] = 16'hffff;
  rom[14302] = 16'hffff;
  rom[14303] = 16'hffde;
  rom[14304] = 16'hffff;
  rom[14305] = 16'hffdf;
  rom[14306] = 16'ha4f3;
  rom[14307] = 16'h2924;
  rom[14308] = 16'h31a6;
  rom[14309] = 16'h9472;
  rom[14310] = 16'hf79e;
  rom[14311] = 16'hffde;
  rom[14312] = 16'hffff;
  rom[14313] = 16'hffff;
  rom[14314] = 16'hffff;
  rom[14315] = 16'hffff;
  rom[14316] = 16'hffff;
  rom[14317] = 16'hffdf;
  rom[14318] = 16'hffdf;
  rom[14319] = 16'hffff;
  rom[14320] = 16'hffff;
  rom[14321] = 16'hffff;
  rom[14322] = 16'hffff;
  rom[14323] = 16'hffff;
  rom[14324] = 16'hffff;
  rom[14325] = 16'hffff;
  rom[14326] = 16'hffff;
  rom[14327] = 16'hffff;
  rom[14328] = 16'hffff;
  rom[14329] = 16'hffff;
  rom[14330] = 16'hffff;
  rom[14331] = 16'hffff;
  rom[14332] = 16'hffff;
  rom[14333] = 16'hffff;
  rom[14334] = 16'hffff;
  rom[14335] = 16'hffff;
  rom[14336] = 16'hffff;
  rom[14337] = 16'hffff;
  rom[14338] = 16'hffff;
  rom[14339] = 16'hffff;
  rom[14340] = 16'hffbe;
  rom[14341] = 16'h8b6b;
  rom[14342] = 16'hc4cb;
  rom[14343] = 16'hf589;
  rom[14344] = 16'hfd49;
  rom[14345] = 16'hf548;
  rom[14346] = 16'hf548;
  rom[14347] = 16'hf528;
  rom[14348] = 16'hfd4a;
  rom[14349] = 16'hfd29;
  rom[14350] = 16'hfd49;
  rom[14351] = 16'hfd27;
  rom[14352] = 16'hf54a;
  rom[14353] = 16'hdd2b;
  rom[14354] = 16'h8347;
  rom[14355] = 16'hde78;
  rom[14356] = 16'hffff;
  rom[14357] = 16'hffff;
  rom[14358] = 16'hffff;
  rom[14359] = 16'hffff;
  rom[14360] = 16'hffff;
  rom[14361] = 16'hffff;
  rom[14362] = 16'hffff;
  rom[14363] = 16'hffff;
  rom[14364] = 16'hffff;
  rom[14365] = 16'hffff;
  rom[14366] = 16'hffff;
  rom[14367] = 16'hffff;
  rom[14368] = 16'hffff;
  rom[14369] = 16'hffff;
  rom[14370] = 16'hffff;
  rom[14371] = 16'hffff;
  rom[14372] = 16'hffff;
  rom[14373] = 16'hffff;
  rom[14374] = 16'hffff;
  rom[14375] = 16'hffff;
  rom[14376] = 16'hffff;
  rom[14377] = 16'hffff;
  rom[14378] = 16'hffff;
  rom[14379] = 16'hffff;
  rom[14380] = 16'hffff;
  rom[14381] = 16'hffff;
  rom[14382] = 16'hffff;
  rom[14383] = 16'hffff;
  rom[14384] = 16'hffff;
  rom[14385] = 16'hffff;
  rom[14386] = 16'hffff;
  rom[14387] = 16'hffff;
  rom[14388] = 16'hffff;
  rom[14389] = 16'hffff;
  rom[14390] = 16'hffff;
  rom[14391] = 16'hffff;
  rom[14392] = 16'hffff;
  rom[14393] = 16'hffff;
  rom[14394] = 16'hffff;
  rom[14395] = 16'hffff;
  rom[14396] = 16'hffff;
  rom[14397] = 16'hffff;
  rom[14398] = 16'hffff;
  rom[14399] = 16'hffff;
  rom[14400] = 16'hffff;
  rom[14401] = 16'hffff;
  rom[14402] = 16'hffff;
  rom[14403] = 16'hffff;
  rom[14404] = 16'hffff;
  rom[14405] = 16'hffff;
  rom[14406] = 16'hffff;
  rom[14407] = 16'hffff;
  rom[14408] = 16'hffff;
  rom[14409] = 16'hffff;
  rom[14410] = 16'hffff;
  rom[14411] = 16'hffff;
  rom[14412] = 16'hffff;
  rom[14413] = 16'hffff;
  rom[14414] = 16'hffff;
  rom[14415] = 16'hffff;
  rom[14416] = 16'hffff;
  rom[14417] = 16'hffff;
  rom[14418] = 16'hffff;
  rom[14419] = 16'hffff;
  rom[14420] = 16'hffff;
  rom[14421] = 16'hffff;
  rom[14422] = 16'hffff;
  rom[14423] = 16'hffff;
  rom[14424] = 16'hffff;
  rom[14425] = 16'hffff;
  rom[14426] = 16'hffff;
  rom[14427] = 16'hffff;
  rom[14428] = 16'hffff;
  rom[14429] = 16'hffff;
  rom[14430] = 16'hffff;
  rom[14431] = 16'hffff;
  rom[14432] = 16'hffff;
  rom[14433] = 16'hffff;
  rom[14434] = 16'hffff;
  rom[14435] = 16'hffff;
  rom[14436] = 16'hffdf;
  rom[14437] = 16'hffff;
  rom[14438] = 16'hffdf;
  rom[14439] = 16'hffdd;
  rom[14440] = 16'ha4ce;
  rom[14441] = 16'hac29;
  rom[14442] = 16'hed4b;
  rom[14443] = 16'hf4e8;
  rom[14444] = 16'hfd28;
  rom[14445] = 16'hfd69;
  rom[14446] = 16'hfd49;
  rom[14447] = 16'hfd68;
  rom[14448] = 16'hf548;
  rom[14449] = 16'hf527;
  rom[14450] = 16'hf568;
  rom[14451] = 16'hed8a;
  rom[14452] = 16'h5a44;
  rom[14453] = 16'hd659;
  rom[14454] = 16'hffdf;
  rom[14455] = 16'hffff;
  rom[14456] = 16'hffff;
  rom[14457] = 16'hffff;
  rom[14458] = 16'hffff;
  rom[14459] = 16'hffff;
  rom[14460] = 16'hffff;
  rom[14461] = 16'hffff;
  rom[14462] = 16'hffff;
  rom[14463] = 16'hffff;
  rom[14464] = 16'hffff;
  rom[14465] = 16'hffff;
  rom[14466] = 16'hffff;
  rom[14467] = 16'hffff;
  rom[14468] = 16'hffff;
  rom[14469] = 16'hffdf;
  rom[14470] = 16'hffff;
  rom[14471] = 16'hffff;
  rom[14472] = 16'hffff;
  rom[14473] = 16'hffff;
  rom[14474] = 16'hff9e;
  rom[14475] = 16'hef5d;
  rom[14476] = 16'hce79;
  rom[14477] = 16'hbdd7;
  rom[14478] = 16'hb595;
  rom[14479] = 16'hbd96;
  rom[14480] = 16'hb5b6;
  rom[14481] = 16'hd658;
  rom[14482] = 16'hef5d;
  rom[14483] = 16'hffbe;
  rom[14484] = 16'hffff;
  rom[14485] = 16'hef3c;
  rom[14486] = 16'h8c50;
  rom[14487] = 16'h5289;
  rom[14488] = 16'he71b;
  rom[14489] = 16'hffff;
  rom[14490] = 16'hffff;
  rom[14491] = 16'hffff;
  rom[14492] = 16'hffff;
  rom[14493] = 16'hffff;
  rom[14494] = 16'hffff;
  rom[14495] = 16'hffff;
  rom[14496] = 16'hffff;
  rom[14497] = 16'hffff;
  rom[14498] = 16'hffff;
  rom[14499] = 16'hffff;
  rom[14500] = 16'hffff;
  rom[14501] = 16'hffff;
  rom[14502] = 16'hffff;
  rom[14503] = 16'hffff;
  rom[14504] = 16'hffff;
  rom[14505] = 16'hf7be;
  rom[14506] = 16'h9492;
  rom[14507] = 16'h4a49;
  rom[14508] = 16'hbdf7;
  rom[14509] = 16'hffff;
  rom[14510] = 16'hffbe;
  rom[14511] = 16'hf79e;
  rom[14512] = 16'he6fb;
  rom[14513] = 16'hc617;
  rom[14514] = 16'had95;
  rom[14515] = 16'had55;
  rom[14516] = 16'hb5b6;
  rom[14517] = 16'hce18;
  rom[14518] = 16'hdeda;
  rom[14519] = 16'hffbe;
  rom[14520] = 16'hffdf;
  rom[14521] = 16'hffff;
  rom[14522] = 16'hffdf;
  rom[14523] = 16'hffff;
  rom[14524] = 16'hffff;
  rom[14525] = 16'hffff;
  rom[14526] = 16'hffff;
  rom[14527] = 16'hffff;
  rom[14528] = 16'hffff;
  rom[14529] = 16'hffff;
  rom[14530] = 16'hffff;
  rom[14531] = 16'hffff;
  rom[14532] = 16'hffff;
  rom[14533] = 16'hffff;
  rom[14534] = 16'hffff;
  rom[14535] = 16'hffff;
  rom[14536] = 16'hffff;
  rom[14537] = 16'hffff;
  rom[14538] = 16'hffdf;
  rom[14539] = 16'hffff;
  rom[14540] = 16'hffff;
  rom[14541] = 16'ha46f;
  rom[14542] = 16'hb469;
  rom[14543] = 16'hf5aa;
  rom[14544] = 16'hf549;
  rom[14545] = 16'hfd68;
  rom[14546] = 16'hfd48;
  rom[14547] = 16'hfd48;
  rom[14548] = 16'hf529;
  rom[14549] = 16'hfd29;
  rom[14550] = 16'hfd07;
  rom[14551] = 16'hfd28;
  rom[14552] = 16'hed49;
  rom[14553] = 16'hd52b;
  rom[14554] = 16'h8ba9;
  rom[14555] = 16'heefa;
  rom[14556] = 16'hffff;
  rom[14557] = 16'hffff;
  rom[14558] = 16'hffff;
  rom[14559] = 16'hffff;
  rom[14560] = 16'hffff;
  rom[14561] = 16'hffff;
  rom[14562] = 16'hffff;
  rom[14563] = 16'hffff;
  rom[14564] = 16'hffff;
  rom[14565] = 16'hffff;
  rom[14566] = 16'hffff;
  rom[14567] = 16'hffff;
  rom[14568] = 16'hffff;
  rom[14569] = 16'hffff;
  rom[14570] = 16'hffff;
  rom[14571] = 16'hffff;
  rom[14572] = 16'hffff;
  rom[14573] = 16'hffff;
  rom[14574] = 16'hffff;
  rom[14575] = 16'hffff;
  rom[14576] = 16'hffff;
  rom[14577] = 16'hffff;
  rom[14578] = 16'hffff;
  rom[14579] = 16'hffff;
  rom[14580] = 16'hffff;
  rom[14581] = 16'hffff;
  rom[14582] = 16'hffff;
  rom[14583] = 16'hffff;
  rom[14584] = 16'hffff;
  rom[14585] = 16'hffff;
  rom[14586] = 16'hffff;
  rom[14587] = 16'hffff;
  rom[14588] = 16'hffff;
  rom[14589] = 16'hffff;
  rom[14590] = 16'hffff;
  rom[14591] = 16'hffff;
  rom[14592] = 16'hffff;
  rom[14593] = 16'hffff;
  rom[14594] = 16'hffff;
  rom[14595] = 16'hffff;
  rom[14596] = 16'hffff;
  rom[14597] = 16'hffff;
  rom[14598] = 16'hffff;
  rom[14599] = 16'hffff;
  rom[14600] = 16'hffff;
  rom[14601] = 16'hffff;
  rom[14602] = 16'hffff;
  rom[14603] = 16'hffff;
  rom[14604] = 16'hffff;
  rom[14605] = 16'hffff;
  rom[14606] = 16'hffff;
  rom[14607] = 16'hffff;
  rom[14608] = 16'hffff;
  rom[14609] = 16'hffff;
  rom[14610] = 16'hffff;
  rom[14611] = 16'hffff;
  rom[14612] = 16'hffff;
  rom[14613] = 16'hffff;
  rom[14614] = 16'hffff;
  rom[14615] = 16'hffff;
  rom[14616] = 16'hffff;
  rom[14617] = 16'hffff;
  rom[14618] = 16'hffff;
  rom[14619] = 16'hffff;
  rom[14620] = 16'hffff;
  rom[14621] = 16'hffff;
  rom[14622] = 16'hffff;
  rom[14623] = 16'hffff;
  rom[14624] = 16'hffff;
  rom[14625] = 16'hffff;
  rom[14626] = 16'hffff;
  rom[14627] = 16'hffff;
  rom[14628] = 16'hffff;
  rom[14629] = 16'hffff;
  rom[14630] = 16'hffff;
  rom[14631] = 16'hffff;
  rom[14632] = 16'hffff;
  rom[14633] = 16'hffff;
  rom[14634] = 16'hffff;
  rom[14635] = 16'hffff;
  rom[14636] = 16'hffff;
  rom[14637] = 16'hffdf;
  rom[14638] = 16'hffff;
  rom[14639] = 16'hffbc;
  rom[14640] = 16'h8389;
  rom[14641] = 16'hbcaa;
  rom[14642] = 16'hed6c;
  rom[14643] = 16'hf54a;
  rom[14644] = 16'hfd4b;
  rom[14645] = 16'hfd4b;
  rom[14646] = 16'hfd09;
  rom[14647] = 16'hfd49;
  rom[14648] = 16'hfd48;
  rom[14649] = 16'hfd48;
  rom[14650] = 16'hfd8a;
  rom[14651] = 16'he54a;
  rom[14652] = 16'h49c2;
  rom[14653] = 16'hef3c;
  rom[14654] = 16'hffff;
  rom[14655] = 16'hffff;
  rom[14656] = 16'hffff;
  rom[14657] = 16'hffff;
  rom[14658] = 16'hffff;
  rom[14659] = 16'hffff;
  rom[14660] = 16'hffff;
  rom[14661] = 16'hffff;
  rom[14662] = 16'hffff;
  rom[14663] = 16'hffff;
  rom[14664] = 16'hffff;
  rom[14665] = 16'hffff;
  rom[14666] = 16'hffff;
  rom[14667] = 16'hffff;
  rom[14668] = 16'hffff;
  rom[14669] = 16'hffff;
  rom[14670] = 16'hffff;
  rom[14671] = 16'hffff;
  rom[14672] = 16'hffdf;
  rom[14673] = 16'hce38;
  rom[14674] = 16'h9472;
  rom[14675] = 16'h528a;
  rom[14676] = 16'h39e6;
  rom[14677] = 16'h1903;
  rom[14678] = 16'h18e3;
  rom[14679] = 16'h2104;
  rom[14680] = 16'h2965;
  rom[14681] = 16'h39c6;
  rom[14682] = 16'h5aaa;
  rom[14683] = 16'h8410;
  rom[14684] = 16'hdebb;
  rom[14685] = 16'hffbe;
  rom[14686] = 16'hf79e;
  rom[14687] = 16'hdedb;
  rom[14688] = 16'hffdf;
  rom[14689] = 16'hffff;
  rom[14690] = 16'hffff;
  rom[14691] = 16'hffff;
  rom[14692] = 16'hffff;
  rom[14693] = 16'hffff;
  rom[14694] = 16'hffff;
  rom[14695] = 16'hffff;
  rom[14696] = 16'hffff;
  rom[14697] = 16'hffff;
  rom[14698] = 16'hffff;
  rom[14699] = 16'hffff;
  rom[14700] = 16'hffff;
  rom[14701] = 16'hffff;
  rom[14702] = 16'hffff;
  rom[14703] = 16'hffff;
  rom[14704] = 16'hffff;
  rom[14705] = 16'hf7de;
  rom[14706] = 16'hef3d;
  rom[14707] = 16'hdedb;
  rom[14708] = 16'hffff;
  rom[14709] = 16'hef7d;
  rom[14710] = 16'hc5d7;
  rom[14711] = 16'h6b4d;
  rom[14712] = 16'h4228;
  rom[14713] = 16'h3185;
  rom[14714] = 16'h2944;
  rom[14715] = 16'h2124;
  rom[14716] = 16'h2103;
  rom[14717] = 16'h2124;
  rom[14718] = 16'h4a28;
  rom[14719] = 16'h6b4c;
  rom[14720] = 16'hb595;
  rom[14721] = 16'hef3c;
  rom[14722] = 16'hffff;
  rom[14723] = 16'hffff;
  rom[14724] = 16'hffff;
  rom[14725] = 16'hffff;
  rom[14726] = 16'hffff;
  rom[14727] = 16'hffff;
  rom[14728] = 16'hffff;
  rom[14729] = 16'hffff;
  rom[14730] = 16'hffff;
  rom[14731] = 16'hffff;
  rom[14732] = 16'hffff;
  rom[14733] = 16'hffff;
  rom[14734] = 16'hffff;
  rom[14735] = 16'hffff;
  rom[14736] = 16'hffff;
  rom[14737] = 16'hffff;
  rom[14738] = 16'hffff;
  rom[14739] = 16'hffff;
  rom[14740] = 16'hffff;
  rom[14741] = 16'hb4f1;
  rom[14742] = 16'hbc8b;
  rom[14743] = 16'hed6a;
  rom[14744] = 16'hf569;
  rom[14745] = 16'hf568;
  rom[14746] = 16'hfd68;
  rom[14747] = 16'hfd68;
  rom[14748] = 16'hfd29;
  rom[14749] = 16'hfd28;
  rom[14750] = 16'hfd28;
  rom[14751] = 16'hfd28;
  rom[14752] = 16'hf54a;
  rom[14753] = 16'hc4cb;
  rom[14754] = 16'h8bcb;
  rom[14755] = 16'hf75b;
  rom[14756] = 16'hffff;
  rom[14757] = 16'hffff;
  rom[14758] = 16'hffff;
  rom[14759] = 16'hffff;
  rom[14760] = 16'hffff;
  rom[14761] = 16'hffff;
  rom[14762] = 16'hffff;
  rom[14763] = 16'hffff;
  rom[14764] = 16'hffff;
  rom[14765] = 16'hffff;
  rom[14766] = 16'hffff;
  rom[14767] = 16'hffff;
  rom[14768] = 16'hffff;
  rom[14769] = 16'hffff;
  rom[14770] = 16'hffff;
  rom[14771] = 16'hffff;
  rom[14772] = 16'hffff;
  rom[14773] = 16'hffff;
  rom[14774] = 16'hffff;
  rom[14775] = 16'hffff;
  rom[14776] = 16'hffff;
  rom[14777] = 16'hffff;
  rom[14778] = 16'hffff;
  rom[14779] = 16'hffff;
  rom[14780] = 16'hffff;
  rom[14781] = 16'hffff;
  rom[14782] = 16'hffff;
  rom[14783] = 16'hffff;
  rom[14784] = 16'hffff;
  rom[14785] = 16'hffff;
  rom[14786] = 16'hffff;
  rom[14787] = 16'hffff;
  rom[14788] = 16'hffff;
  rom[14789] = 16'hffff;
  rom[14790] = 16'hffff;
  rom[14791] = 16'hffff;
  rom[14792] = 16'hffff;
  rom[14793] = 16'hffff;
  rom[14794] = 16'hffff;
  rom[14795] = 16'hffff;
  rom[14796] = 16'hffff;
  rom[14797] = 16'hffff;
  rom[14798] = 16'hffff;
  rom[14799] = 16'hffff;
  rom[14800] = 16'hffff;
  rom[14801] = 16'hffff;
  rom[14802] = 16'hffff;
  rom[14803] = 16'hffff;
  rom[14804] = 16'hffff;
  rom[14805] = 16'hffff;
  rom[14806] = 16'hffff;
  rom[14807] = 16'hffff;
  rom[14808] = 16'hffff;
  rom[14809] = 16'hffff;
  rom[14810] = 16'hffff;
  rom[14811] = 16'hffff;
  rom[14812] = 16'hffff;
  rom[14813] = 16'hffff;
  rom[14814] = 16'hffff;
  rom[14815] = 16'hffff;
  rom[14816] = 16'hffff;
  rom[14817] = 16'hffff;
  rom[14818] = 16'hffff;
  rom[14819] = 16'hffff;
  rom[14820] = 16'hffff;
  rom[14821] = 16'hffff;
  rom[14822] = 16'hffff;
  rom[14823] = 16'hffff;
  rom[14824] = 16'hffff;
  rom[14825] = 16'hffff;
  rom[14826] = 16'hffff;
  rom[14827] = 16'hffff;
  rom[14828] = 16'hffff;
  rom[14829] = 16'hffff;
  rom[14830] = 16'hffff;
  rom[14831] = 16'hffff;
  rom[14832] = 16'hffdf;
  rom[14833] = 16'hffff;
  rom[14834] = 16'hffff;
  rom[14835] = 16'hffff;
  rom[14836] = 16'hffde;
  rom[14837] = 16'hff9d;
  rom[14838] = 16'hffbc;
  rom[14839] = 16'hde96;
  rom[14840] = 16'h6283;
  rom[14841] = 16'hb469;
  rom[14842] = 16'hdd4b;
  rom[14843] = 16'he52a;
  rom[14844] = 16'hed0b;
  rom[14845] = 16'hfd8d;
  rom[14846] = 16'hf52a;
  rom[14847] = 16'hf528;
  rom[14848] = 16'hfd28;
  rom[14849] = 16'hfd49;
  rom[14850] = 16'hf56a;
  rom[14851] = 16'hdd0a;
  rom[14852] = 16'h51e2;
  rom[14853] = 16'hff9d;
  rom[14854] = 16'hffff;
  rom[14855] = 16'hffff;
  rom[14856] = 16'hffff;
  rom[14857] = 16'hffff;
  rom[14858] = 16'hffff;
  rom[14859] = 16'hffff;
  rom[14860] = 16'hffff;
  rom[14861] = 16'hffff;
  rom[14862] = 16'hffff;
  rom[14863] = 16'hffff;
  rom[14864] = 16'hffff;
  rom[14865] = 16'hffff;
  rom[14866] = 16'hffff;
  rom[14867] = 16'hffff;
  rom[14868] = 16'hffff;
  rom[14869] = 16'hffff;
  rom[14870] = 16'hffdf;
  rom[14871] = 16'hef3c;
  rom[14872] = 16'h9c92;
  rom[14873] = 16'h4a28;
  rom[14874] = 16'h0861;
  rom[14875] = 16'h18e3;
  rom[14876] = 16'h1081;
  rom[14877] = 16'h2103;
  rom[14878] = 16'h18e2;
  rom[14879] = 16'h1081;
  rom[14880] = 16'h10a1;
  rom[14881] = 16'h1081;
  rom[14882] = 16'h2103;
  rom[14883] = 16'h18e3;
  rom[14884] = 16'h2965;
  rom[14885] = 16'ha514;
  rom[14886] = 16'hf77d;
  rom[14887] = 16'hffff;
  rom[14888] = 16'hffff;
  rom[14889] = 16'hffff;
  rom[14890] = 16'hffff;
  rom[14891] = 16'hffff;
  rom[14892] = 16'hffff;
  rom[14893] = 16'hffff;
  rom[14894] = 16'hffff;
  rom[14895] = 16'hffff;
  rom[14896] = 16'hffff;
  rom[14897] = 16'hffff;
  rom[14898] = 16'hffff;
  rom[14899] = 16'hffff;
  rom[14900] = 16'hffff;
  rom[14901] = 16'hffff;
  rom[14902] = 16'hffff;
  rom[14903] = 16'hffdf;
  rom[14904] = 16'hffdf;
  rom[14905] = 16'hffff;
  rom[14906] = 16'hffff;
  rom[14907] = 16'hffdf;
  rom[14908] = 16'hc638;
  rom[14909] = 16'h6b4d;
  rom[14910] = 16'h18e2;
  rom[14911] = 16'h2124;
  rom[14912] = 16'h10a2;
  rom[14913] = 16'h18a2;
  rom[14914] = 16'h1081;
  rom[14915] = 16'h10a1;
  rom[14916] = 16'h1903;
  rom[14917] = 16'h2103;
  rom[14918] = 16'h10a1;
  rom[14919] = 16'h10a1;
  rom[14920] = 16'h1903;
  rom[14921] = 16'h7bae;
  rom[14922] = 16'hc617;
  rom[14923] = 16'hffbf;
  rom[14924] = 16'hffff;
  rom[14925] = 16'hffff;
  rom[14926] = 16'hffff;
  rom[14927] = 16'hffff;
  rom[14928] = 16'hffff;
  rom[14929] = 16'hffff;
  rom[14930] = 16'hffff;
  rom[14931] = 16'hffff;
  rom[14932] = 16'hffff;
  rom[14933] = 16'hffff;
  rom[14934] = 16'hffff;
  rom[14935] = 16'hffff;
  rom[14936] = 16'hffff;
  rom[14937] = 16'hffff;
  rom[14938] = 16'hffff;
  rom[14939] = 16'hffff;
  rom[14940] = 16'hffff;
  rom[14941] = 16'hc554;
  rom[14942] = 16'hac29;
  rom[14943] = 16'hed6a;
  rom[14944] = 16'hf569;
  rom[14945] = 16'hfd68;
  rom[14946] = 16'hf547;
  rom[14947] = 16'hfd89;
  rom[14948] = 16'hfd28;
  rom[14949] = 16'hfd29;
  rom[14950] = 16'hfd08;
  rom[14951] = 16'hfd48;
  rom[14952] = 16'hed2a;
  rom[14953] = 16'hb469;
  rom[14954] = 16'h93eb;
  rom[14955] = 16'hff9d;
  rom[14956] = 16'hffff;
  rom[14957] = 16'hffdf;
  rom[14958] = 16'hffff;
  rom[14959] = 16'hffff;
  rom[14960] = 16'hffff;
  rom[14961] = 16'hffff;
  rom[14962] = 16'hffff;
  rom[14963] = 16'hffff;
  rom[14964] = 16'hffff;
  rom[14965] = 16'hffff;
  rom[14966] = 16'hffff;
  rom[14967] = 16'hffff;
  rom[14968] = 16'hffff;
  rom[14969] = 16'hffff;
  rom[14970] = 16'hffff;
  rom[14971] = 16'hffff;
  rom[14972] = 16'hffff;
  rom[14973] = 16'hffff;
  rom[14974] = 16'hffff;
  rom[14975] = 16'hffff;
  rom[14976] = 16'hffff;
  rom[14977] = 16'hffff;
  rom[14978] = 16'hffff;
  rom[14979] = 16'hffff;
  rom[14980] = 16'hffff;
  rom[14981] = 16'hffff;
  rom[14982] = 16'hffff;
  rom[14983] = 16'hffff;
  rom[14984] = 16'hffff;
  rom[14985] = 16'hffff;
  rom[14986] = 16'hffff;
  rom[14987] = 16'hffff;
  rom[14988] = 16'hffff;
  rom[14989] = 16'hffff;
  rom[14990] = 16'hffff;
  rom[14991] = 16'hffff;
  rom[14992] = 16'hffff;
  rom[14993] = 16'hffff;
  rom[14994] = 16'hffff;
  rom[14995] = 16'hffff;
  rom[14996] = 16'hffff;
  rom[14997] = 16'hffff;
  rom[14998] = 16'hffff;
  rom[14999] = 16'hffff;
  rom[15000] = 16'hffff;
  rom[15001] = 16'hffff;
  rom[15002] = 16'hffff;
  rom[15003] = 16'hffff;
  rom[15004] = 16'hffff;
  rom[15005] = 16'hffff;
  rom[15006] = 16'hffff;
  rom[15007] = 16'hffff;
  rom[15008] = 16'hffff;
  rom[15009] = 16'hffff;
  rom[15010] = 16'hffff;
  rom[15011] = 16'hffff;
  rom[15012] = 16'hffff;
  rom[15013] = 16'hffff;
  rom[15014] = 16'hffff;
  rom[15015] = 16'hffff;
  rom[15016] = 16'hffff;
  rom[15017] = 16'hffff;
  rom[15018] = 16'hffff;
  rom[15019] = 16'hffff;
  rom[15020] = 16'hffff;
  rom[15021] = 16'hffff;
  rom[15022] = 16'hffff;
  rom[15023] = 16'hffff;
  rom[15024] = 16'hffff;
  rom[15025] = 16'hffff;
  rom[15026] = 16'hffff;
  rom[15027] = 16'hffff;
  rom[15028] = 16'hffff;
  rom[15029] = 16'hffdf;
  rom[15030] = 16'hffff;
  rom[15031] = 16'hffff;
  rom[15032] = 16'hffff;
  rom[15033] = 16'hffdd;
  rom[15034] = 16'hef1a;
  rom[15035] = 16'hb572;
  rom[15036] = 16'h9c6d;
  rom[15037] = 16'h7bc9;
  rom[15038] = 16'h8c0a;
  rom[15039] = 16'h6b26;
  rom[15040] = 16'h6ac3;
  rom[15041] = 16'h8302;
  rom[15042] = 16'h82a2;
  rom[15043] = 16'h8ae2;
  rom[15044] = 16'ha344;
  rom[15045] = 16'hc448;
  rom[15046] = 16'hf56c;
  rom[15047] = 16'hf549;
  rom[15048] = 16'hfd49;
  rom[15049] = 16'hfd29;
  rom[15050] = 16'hfd6b;
  rom[15051] = 16'hdce9;
  rom[15052] = 16'h6264;
  rom[15053] = 16'hffdd;
  rom[15054] = 16'hffff;
  rom[15055] = 16'hffff;
  rom[15056] = 16'hffff;
  rom[15057] = 16'hffff;
  rom[15058] = 16'hffff;
  rom[15059] = 16'hffff;
  rom[15060] = 16'hffff;
  rom[15061] = 16'hffff;
  rom[15062] = 16'hffff;
  rom[15063] = 16'hffff;
  rom[15064] = 16'hffff;
  rom[15065] = 16'hffff;
  rom[15066] = 16'hffff;
  rom[15067] = 16'hffff;
  rom[15068] = 16'hffff;
  rom[15069] = 16'hffdf;
  rom[15070] = 16'hdedb;
  rom[15071] = 16'h738d;
  rom[15072] = 16'h2944;
  rom[15073] = 16'h1061;
  rom[15074] = 16'h2104;
  rom[15075] = 16'h10a2;
  rom[15076] = 16'h20e3;
  rom[15077] = 16'h10a2;
  rom[15078] = 16'h10c2;
  rom[15079] = 16'h10a2;
  rom[15080] = 16'h20c2;
  rom[15081] = 16'h18a2;
  rom[15082] = 16'h18c3;
  rom[15083] = 16'h18c2;
  rom[15084] = 16'h20c3;
  rom[15085] = 16'h2924;
  rom[15086] = 16'h7b8d;
  rom[15087] = 16'hdedb;
  rom[15088] = 16'hffff;
  rom[15089] = 16'hffff;
  rom[15090] = 16'hffff;
  rom[15091] = 16'hffff;
  rom[15092] = 16'hffff;
  rom[15093] = 16'hffff;
  rom[15094] = 16'hffff;
  rom[15095] = 16'hffff;
  rom[15096] = 16'hffff;
  rom[15097] = 16'hffff;
  rom[15098] = 16'hffff;
  rom[15099] = 16'hffff;
  rom[15100] = 16'hffff;
  rom[15101] = 16'hffff;
  rom[15102] = 16'hffff;
  rom[15103] = 16'hffdf;
  rom[15104] = 16'hffff;
  rom[15105] = 16'hffff;
  rom[15106] = 16'hffdf;
  rom[15107] = 16'hb596;
  rom[15108] = 16'h5269;
  rom[15109] = 16'h18c2;
  rom[15110] = 16'h18c3;
  rom[15111] = 16'h10a2;
  rom[15112] = 16'h18c3;
  rom[15113] = 16'h18c2;
  rom[15114] = 16'h20e3;
  rom[15115] = 16'h10a2;
  rom[15116] = 16'h18a2;
  rom[15117] = 16'h18c2;
  rom[15118] = 16'h18c2;
  rom[15119] = 16'h18c2;
  rom[15120] = 16'h18a3;
  rom[15121] = 16'h18a2;
  rom[15122] = 16'h4228;
  rom[15123] = 16'had34;
  rom[15124] = 16'hffbf;
  rom[15125] = 16'hffff;
  rom[15126] = 16'hffff;
  rom[15127] = 16'hffff;
  rom[15128] = 16'hffff;
  rom[15129] = 16'hffff;
  rom[15130] = 16'hffff;
  rom[15131] = 16'hffff;
  rom[15132] = 16'hffff;
  rom[15133] = 16'hffff;
  rom[15134] = 16'hffff;
  rom[15135] = 16'hffff;
  rom[15136] = 16'hffff;
  rom[15137] = 16'hffff;
  rom[15138] = 16'hffff;
  rom[15139] = 16'hffff;
  rom[15140] = 16'hffff;
  rom[15141] = 16'hc554;
  rom[15142] = 16'hb44a;
  rom[15143] = 16'hed6a;
  rom[15144] = 16'hf569;
  rom[15145] = 16'hfd68;
  rom[15146] = 16'hfd47;
  rom[15147] = 16'hfd68;
  rom[15148] = 16'hfd49;
  rom[15149] = 16'hfd29;
  rom[15150] = 16'hfd4a;
  rom[15151] = 16'hfd48;
  rom[15152] = 16'hed4a;
  rom[15153] = 16'habe9;
  rom[15154] = 16'hb4f1;
  rom[15155] = 16'hfffe;
  rom[15156] = 16'hffff;
  rom[15157] = 16'hffff;
  rom[15158] = 16'hffff;
  rom[15159] = 16'hffff;
  rom[15160] = 16'hffff;
  rom[15161] = 16'hffff;
  rom[15162] = 16'hffff;
  rom[15163] = 16'hffff;
  rom[15164] = 16'hffff;
  rom[15165] = 16'hffff;
  rom[15166] = 16'hffff;
  rom[15167] = 16'hffff;
  rom[15168] = 16'hffff;
  rom[15169] = 16'hffff;
  rom[15170] = 16'hffff;
  rom[15171] = 16'hffff;
  rom[15172] = 16'hffff;
  rom[15173] = 16'hffff;
  rom[15174] = 16'hffff;
  rom[15175] = 16'hffff;
  rom[15176] = 16'hffff;
  rom[15177] = 16'hffff;
  rom[15178] = 16'hffff;
  rom[15179] = 16'hffff;
  rom[15180] = 16'hffff;
  rom[15181] = 16'hffff;
  rom[15182] = 16'hffff;
  rom[15183] = 16'hffff;
  rom[15184] = 16'hffff;
  rom[15185] = 16'hffff;
  rom[15186] = 16'hffff;
  rom[15187] = 16'hffff;
  rom[15188] = 16'hffff;
  rom[15189] = 16'hffff;
  rom[15190] = 16'hffff;
  rom[15191] = 16'hffff;
  rom[15192] = 16'hffff;
  rom[15193] = 16'hffff;
  rom[15194] = 16'hffff;
  rom[15195] = 16'hffff;
  rom[15196] = 16'hffff;
  rom[15197] = 16'hffff;
  rom[15198] = 16'hffff;
  rom[15199] = 16'hffff;
  rom[15200] = 16'hffff;
  rom[15201] = 16'hffff;
  rom[15202] = 16'hffff;
  rom[15203] = 16'hffff;
  rom[15204] = 16'hffff;
  rom[15205] = 16'hffff;
  rom[15206] = 16'hffff;
  rom[15207] = 16'hffff;
  rom[15208] = 16'hffff;
  rom[15209] = 16'hffff;
  rom[15210] = 16'hffff;
  rom[15211] = 16'hffff;
  rom[15212] = 16'hffff;
  rom[15213] = 16'hffff;
  rom[15214] = 16'hffff;
  rom[15215] = 16'hffff;
  rom[15216] = 16'hffff;
  rom[15217] = 16'hffff;
  rom[15218] = 16'hffff;
  rom[15219] = 16'hffff;
  rom[15220] = 16'hffff;
  rom[15221] = 16'hffff;
  rom[15222] = 16'hffff;
  rom[15223] = 16'hffff;
  rom[15224] = 16'hffff;
  rom[15225] = 16'hffff;
  rom[15226] = 16'hffdf;
  rom[15227] = 16'hffff;
  rom[15228] = 16'hffff;
  rom[15229] = 16'hffff;
  rom[15230] = 16'hff9d;
  rom[15231] = 16'hfffd;
  rom[15232] = 16'hf779;
  rom[15233] = 16'had2f;
  rom[15234] = 16'h6b06;
  rom[15235] = 16'h7b47;
  rom[15236] = 16'h9407;
  rom[15237] = 16'hacea;
  rom[15238] = 16'hc5ec;
  rom[15239] = 16'he68f;
  rom[15240] = 16'he68e;
  rom[15241] = 16'hddeb;
  rom[15242] = 16'hcd48;
  rom[15243] = 16'hbca7;
  rom[15244] = 16'h8342;
  rom[15245] = 16'h7260;
  rom[15246] = 16'h8b03;
  rom[15247] = 16'hed6a;
  rom[15248] = 16'hf569;
  rom[15249] = 16'hfd29;
  rom[15250] = 16'hfd6a;
  rom[15251] = 16'hdd2a;
  rom[15252] = 16'h49e2;
  rom[15253] = 16'hffdd;
  rom[15254] = 16'hffff;
  rom[15255] = 16'hffff;
  rom[15256] = 16'hffff;
  rom[15257] = 16'hffff;
  rom[15258] = 16'hffff;
  rom[15259] = 16'hffff;
  rom[15260] = 16'hffff;
  rom[15261] = 16'hffff;
  rom[15262] = 16'hffff;
  rom[15263] = 16'hffff;
  rom[15264] = 16'hffdf;
  rom[15265] = 16'hffff;
  rom[15266] = 16'hffdf;
  rom[15267] = 16'hffff;
  rom[15268] = 16'hffde;
  rom[15269] = 16'hffbe;
  rom[15270] = 16'h6b6d;
  rom[15271] = 16'h18e3;
  rom[15272] = 16'h18c2;
  rom[15273] = 16'h18c2;
  rom[15274] = 16'h1061;
  rom[15275] = 16'h18c3;
  rom[15276] = 16'h1081;
  rom[15277] = 16'h18e3;
  rom[15278] = 16'h18c2;
  rom[15279] = 16'h18c2;
  rom[15280] = 16'h10c2;
  rom[15281] = 16'h18c2;
  rom[15282] = 16'h1081;
  rom[15283] = 16'h18e3;
  rom[15284] = 16'h10a2;
  rom[15285] = 16'h10a2;
  rom[15286] = 16'h2123;
  rom[15287] = 16'h6b4d;
  rom[15288] = 16'hf79e;
  rom[15289] = 16'hffff;
  rom[15290] = 16'hffff;
  rom[15291] = 16'hffff;
  rom[15292] = 16'hffff;
  rom[15293] = 16'hffff;
  rom[15294] = 16'hffff;
  rom[15295] = 16'hffff;
  rom[15296] = 16'hffff;
  rom[15297] = 16'hffff;
  rom[15298] = 16'hffff;
  rom[15299] = 16'hffff;
  rom[15300] = 16'hffff;
  rom[15301] = 16'hffff;
  rom[15302] = 16'hffff;
  rom[15303] = 16'hffff;
  rom[15304] = 16'hffde;
  rom[15305] = 16'hffff;
  rom[15306] = 16'hb596;
  rom[15307] = 16'h4228;
  rom[15308] = 16'h1081;
  rom[15309] = 16'h20e3;
  rom[15310] = 16'h18a2;
  rom[15311] = 16'h18a2;
  rom[15312] = 16'h18c2;
  rom[15313] = 16'h18a2;
  rom[15314] = 16'h1081;
  rom[15315] = 16'h18c2;
  rom[15316] = 16'h18c2;
  rom[15317] = 16'h10c2;
  rom[15318] = 16'h10c2;
  rom[15319] = 16'h10a2;
  rom[15320] = 16'h10a1;
  rom[15321] = 16'h1061;
  rom[15322] = 16'h2103;
  rom[15323] = 16'h41e7;
  rom[15324] = 16'had35;
  rom[15325] = 16'hffdf;
  rom[15326] = 16'hffff;
  rom[15327] = 16'hffff;
  rom[15328] = 16'hffff;
  rom[15329] = 16'hffff;
  rom[15330] = 16'hffff;
  rom[15331] = 16'hffff;
  rom[15332] = 16'hffff;
  rom[15333] = 16'hffff;
  rom[15334] = 16'hffff;
  rom[15335] = 16'hffff;
  rom[15336] = 16'hffff;
  rom[15337] = 16'hffff;
  rom[15338] = 16'hffff;
  rom[15339] = 16'hffff;
  rom[15340] = 16'hffff;
  rom[15341] = 16'hbd33;
  rom[15342] = 16'hb46a;
  rom[15343] = 16'hed8a;
  rom[15344] = 16'hed48;
  rom[15345] = 16'hfd68;
  rom[15346] = 16'hf527;
  rom[15347] = 16'hfd48;
  rom[15348] = 16'hf528;
  rom[15349] = 16'hfd29;
  rom[15350] = 16'hfd29;
  rom[15351] = 16'hf529;
  rom[15352] = 16'he52a;
  rom[15353] = 16'habe9;
  rom[15354] = 16'hcd94;
  rom[15355] = 16'hffff;
  rom[15356] = 16'hffdf;
  rom[15357] = 16'hffff;
  rom[15358] = 16'hffff;
  rom[15359] = 16'hffff;
  rom[15360] = 16'hffff;
  rom[15361] = 16'hffff;
  rom[15362] = 16'hffff;
  rom[15363] = 16'hffff;
  rom[15364] = 16'hffff;
  rom[15365] = 16'hffff;
  rom[15366] = 16'hffff;
  rom[15367] = 16'hffff;
  rom[15368] = 16'hffff;
  rom[15369] = 16'hffff;
  rom[15370] = 16'hffff;
  rom[15371] = 16'hffff;
  rom[15372] = 16'hffff;
  rom[15373] = 16'hffff;
  rom[15374] = 16'hffff;
  rom[15375] = 16'hffff;
  rom[15376] = 16'hffff;
  rom[15377] = 16'hffff;
  rom[15378] = 16'hffff;
  rom[15379] = 16'hffff;
  rom[15380] = 16'hffff;
  rom[15381] = 16'hffff;
  rom[15382] = 16'hffff;
  rom[15383] = 16'hffff;
  rom[15384] = 16'hffff;
  rom[15385] = 16'hffff;
  rom[15386] = 16'hffff;
  rom[15387] = 16'hffff;
  rom[15388] = 16'hffff;
  rom[15389] = 16'hffff;
  rom[15390] = 16'hffff;
  rom[15391] = 16'hffff;
  rom[15392] = 16'hffff;
  rom[15393] = 16'hffff;
  rom[15394] = 16'hffff;
  rom[15395] = 16'hffff;
  rom[15396] = 16'hffff;
  rom[15397] = 16'hffff;
  rom[15398] = 16'hffff;
  rom[15399] = 16'hffff;
  rom[15400] = 16'hffff;
  rom[15401] = 16'hffff;
  rom[15402] = 16'hffff;
  rom[15403] = 16'hffff;
  rom[15404] = 16'hffff;
  rom[15405] = 16'hffff;
  rom[15406] = 16'hffff;
  rom[15407] = 16'hffff;
  rom[15408] = 16'hffff;
  rom[15409] = 16'hffff;
  rom[15410] = 16'hffff;
  rom[15411] = 16'hffff;
  rom[15412] = 16'hffff;
  rom[15413] = 16'hffff;
  rom[15414] = 16'hffff;
  rom[15415] = 16'hffff;
  rom[15416] = 16'hffff;
  rom[15417] = 16'hffff;
  rom[15418] = 16'hffff;
  rom[15419] = 16'hffff;
  rom[15420] = 16'hffff;
  rom[15421] = 16'hffff;
  rom[15422] = 16'hffff;
  rom[15423] = 16'hffff;
  rom[15424] = 16'hffff;
  rom[15425] = 16'hffff;
  rom[15426] = 16'hffff;
  rom[15427] = 16'hffff;
  rom[15428] = 16'hffff;
  rom[15429] = 16'hffff;
  rom[15430] = 16'hfffe;
  rom[15431] = 16'hded7;
  rom[15432] = 16'h83e9;
  rom[15433] = 16'h6b03;
  rom[15434] = 16'hacea;
  rom[15435] = 16'hde2d;
  rom[15436] = 16'hf6ee;
  rom[15437] = 16'hf70c;
  rom[15438] = 16'hf70c;
  rom[15439] = 16'hf70c;
  rom[15440] = 16'hff2c;
  rom[15441] = 16'hf6eb;
  rom[15442] = 16'hff0c;
  rom[15443] = 16'hf6ec;
  rom[15444] = 16'heecc;
  rom[15445] = 16'hb4e6;
  rom[15446] = 16'h8302;
  rom[15447] = 16'hb3e4;
  rom[15448] = 16'hed4a;
  rom[15449] = 16'hf56a;
  rom[15450] = 16'hf54a;
  rom[15451] = 16'he54a;
  rom[15452] = 16'h51c2;
  rom[15453] = 16'hef5c;
  rom[15454] = 16'hffff;
  rom[15455] = 16'hffff;
  rom[15456] = 16'hffff;
  rom[15457] = 16'hffff;
  rom[15458] = 16'hffff;
  rom[15459] = 16'hffff;
  rom[15460] = 16'hffff;
  rom[15461] = 16'hffff;
  rom[15462] = 16'hffff;
  rom[15463] = 16'hffff;
  rom[15464] = 16'hffff;
  rom[15465] = 16'hffff;
  rom[15466] = 16'hffff;
  rom[15467] = 16'hffff;
  rom[15468] = 16'hffbf;
  rom[15469] = 16'h8410;
  rom[15470] = 16'h2103;
  rom[15471] = 16'h20e3;
  rom[15472] = 16'h1082;
  rom[15473] = 16'h18e2;
  rom[15474] = 16'h20c3;
  rom[15475] = 16'h18a2;
  rom[15476] = 16'h18c2;
  rom[15477] = 16'h10a2;
  rom[15478] = 16'h18c3;
  rom[15479] = 16'h10a2;
  rom[15480] = 16'h18c2;
  rom[15481] = 16'h18c2;
  rom[15482] = 16'h18c2;
  rom[15483] = 16'h18c2;
  rom[15484] = 16'h18c2;
  rom[15485] = 16'h10a2;
  rom[15486] = 16'h18c2;
  rom[15487] = 16'h2123;
  rom[15488] = 16'h9471;
  rom[15489] = 16'hffbe;
  rom[15490] = 16'hffff;
  rom[15491] = 16'hffff;
  rom[15492] = 16'hffff;
  rom[15493] = 16'hffff;
  rom[15494] = 16'hffff;
  rom[15495] = 16'hffff;
  rom[15496] = 16'hffff;
  rom[15497] = 16'hffff;
  rom[15498] = 16'hffff;
  rom[15499] = 16'hffff;
  rom[15500] = 16'hffff;
  rom[15501] = 16'hffff;
  rom[15502] = 16'hffff;
  rom[15503] = 16'hffde;
  rom[15504] = 16'hffff;
  rom[15505] = 16'hdefb;
  rom[15506] = 16'h41e7;
  rom[15507] = 16'h1081;
  rom[15508] = 16'h18e3;
  rom[15509] = 16'h18c2;
  rom[15510] = 16'h18a2;
  rom[15511] = 16'h18e2;
  rom[15512] = 16'h18c2;
  rom[15513] = 16'h18a2;
  rom[15514] = 16'h18c3;
  rom[15515] = 16'h18a2;
  rom[15516] = 16'h18a2;
  rom[15517] = 16'h10c2;
  rom[15518] = 16'h18c2;
  rom[15519] = 16'h18c2;
  rom[15520] = 16'h10c2;
  rom[15521] = 16'h18c2;
  rom[15522] = 16'h18a2;
  rom[15523] = 16'h1061;
  rom[15524] = 16'h4a69;
  rom[15525] = 16'hc618;
  rom[15526] = 16'hffff;
  rom[15527] = 16'hffff;
  rom[15528] = 16'hffff;
  rom[15529] = 16'hffff;
  rom[15530] = 16'hffff;
  rom[15531] = 16'hffff;
  rom[15532] = 16'hffff;
  rom[15533] = 16'hffff;
  rom[15534] = 16'hffff;
  rom[15535] = 16'hffff;
  rom[15536] = 16'hffff;
  rom[15537] = 16'hffff;
  rom[15538] = 16'hffff;
  rom[15539] = 16'hffff;
  rom[15540] = 16'hffff;
  rom[15541] = 16'hbd33;
  rom[15542] = 16'hb44a;
  rom[15543] = 16'hed4a;
  rom[15544] = 16'hf56a;
  rom[15545] = 16'hfd48;
  rom[15546] = 16'hfd68;
  rom[15547] = 16'hfd28;
  rom[15548] = 16'hfd49;
  rom[15549] = 16'hf529;
  rom[15550] = 16'hfd4a;
  rom[15551] = 16'hf529;
  rom[15552] = 16'hed6b;
  rom[15553] = 16'ha3e9;
  rom[15554] = 16'hddf7;
  rom[15555] = 16'hffff;
  rom[15556] = 16'hffff;
  rom[15557] = 16'hffff;
  rom[15558] = 16'hffff;
  rom[15559] = 16'hffff;
  rom[15560] = 16'hffff;
  rom[15561] = 16'hffff;
  rom[15562] = 16'hffff;
  rom[15563] = 16'hffff;
  rom[15564] = 16'hffff;
  rom[15565] = 16'hffff;
  rom[15566] = 16'hffff;
  rom[15567] = 16'hffff;
  rom[15568] = 16'hffff;
  rom[15569] = 16'hffff;
  rom[15570] = 16'hffff;
  rom[15571] = 16'hffff;
  rom[15572] = 16'hffff;
  rom[15573] = 16'hffff;
  rom[15574] = 16'hffff;
  rom[15575] = 16'hffff;
  rom[15576] = 16'hffff;
  rom[15577] = 16'hffff;
  rom[15578] = 16'hffff;
  rom[15579] = 16'hffff;
  rom[15580] = 16'hffff;
  rom[15581] = 16'hffff;
  rom[15582] = 16'hffff;
  rom[15583] = 16'hffff;
  rom[15584] = 16'hffff;
  rom[15585] = 16'hffff;
  rom[15586] = 16'hffff;
  rom[15587] = 16'hffff;
  rom[15588] = 16'hffff;
  rom[15589] = 16'hffff;
  rom[15590] = 16'hffff;
  rom[15591] = 16'hffff;
  rom[15592] = 16'hffff;
  rom[15593] = 16'hffff;
  rom[15594] = 16'hffff;
  rom[15595] = 16'hffff;
  rom[15596] = 16'hffff;
  rom[15597] = 16'hffff;
  rom[15598] = 16'hffff;
  rom[15599] = 16'hffff;
  rom[15600] = 16'hffff;
  rom[15601] = 16'hffff;
  rom[15602] = 16'hffff;
  rom[15603] = 16'hffff;
  rom[15604] = 16'hffff;
  rom[15605] = 16'hffff;
  rom[15606] = 16'hffff;
  rom[15607] = 16'hffff;
  rom[15608] = 16'hffff;
  rom[15609] = 16'hffff;
  rom[15610] = 16'hffff;
  rom[15611] = 16'hffff;
  rom[15612] = 16'hffff;
  rom[15613] = 16'hffff;
  rom[15614] = 16'hffff;
  rom[15615] = 16'hffff;
  rom[15616] = 16'hffff;
  rom[15617] = 16'hffff;
  rom[15618] = 16'hffff;
  rom[15619] = 16'hffff;
  rom[15620] = 16'hffff;
  rom[15621] = 16'hffff;
  rom[15622] = 16'hffff;
  rom[15623] = 16'hffff;
  rom[15624] = 16'hffdf;
  rom[15625] = 16'hffff;
  rom[15626] = 16'hffff;
  rom[15627] = 16'hffff;
  rom[15628] = 16'hffff;
  rom[15629] = 16'hfffe;
  rom[15630] = 16'hce35;
  rom[15631] = 16'h6b06;
  rom[15632] = 16'h83e6;
  rom[15633] = 16'he68f;
  rom[15634] = 16'heecd;
  rom[15635] = 16'hff0c;
  rom[15636] = 16'hf70a;
  rom[15637] = 16'hff4a;
  rom[15638] = 16'hef08;
  rom[15639] = 16'hf74a;
  rom[15640] = 16'hf729;
  rom[15641] = 16'hff4a;
  rom[15642] = 16'hf72a;
  rom[15643] = 16'hf72a;
  rom[15644] = 16'hef2b;
  rom[15645] = 16'he6ab;
  rom[15646] = 16'hb4e6;
  rom[15647] = 16'h7260;
  rom[15648] = 16'hd4e9;
  rom[15649] = 16'hf56b;
  rom[15650] = 16'hed48;
  rom[15651] = 16'he56a;
  rom[15652] = 16'h51e2;
  rom[15653] = 16'he6ba;
  rom[15654] = 16'hffdf;
  rom[15655] = 16'hffff;
  rom[15656] = 16'hffff;
  rom[15657] = 16'hffff;
  rom[15658] = 16'hffff;
  rom[15659] = 16'hffff;
  rom[15660] = 16'hffff;
  rom[15661] = 16'hffff;
  rom[15662] = 16'hffff;
  rom[15663] = 16'hffff;
  rom[15664] = 16'hffff;
  rom[15665] = 16'hffff;
  rom[15666] = 16'hffff;
  rom[15667] = 16'hffff;
  rom[15668] = 16'hbdb6;
  rom[15669] = 16'h3145;
  rom[15670] = 16'h10a2;
  rom[15671] = 16'h18e3;
  rom[15672] = 16'h1082;
  rom[15673] = 16'h20e3;
  rom[15674] = 16'h0840;
  rom[15675] = 16'h20c3;
  rom[15676] = 16'h1082;
  rom[15677] = 16'h18c3;
  rom[15678] = 16'h10a2;
  rom[15679] = 16'h18c2;
  rom[15680] = 16'h10a2;
  rom[15681] = 16'h18c2;
  rom[15682] = 16'h10c2;
  rom[15683] = 16'h10a2;
  rom[15684] = 16'h18c2;
  rom[15685] = 16'h18a2;
  rom[15686] = 16'h18c2;
  rom[15687] = 16'h18a2;
  rom[15688] = 16'h10a1;
  rom[15689] = 16'hce38;
  rom[15690] = 16'hffbe;
  rom[15691] = 16'hffff;
  rom[15692] = 16'hffff;
  rom[15693] = 16'hffff;
  rom[15694] = 16'hffff;
  rom[15695] = 16'hffff;
  rom[15696] = 16'hffff;
  rom[15697] = 16'hffff;
  rom[15698] = 16'hffff;
  rom[15699] = 16'hffff;
  rom[15700] = 16'hffff;
  rom[15701] = 16'hffff;
  rom[15702] = 16'hffff;
  rom[15703] = 16'hffdf;
  rom[15704] = 16'hffff;
  rom[15705] = 16'h62eb;
  rom[15706] = 16'h10c2;
  rom[15707] = 16'h18e3;
  rom[15708] = 16'h10a2;
  rom[15709] = 16'h18a2;
  rom[15710] = 16'h10c2;
  rom[15711] = 16'h18a2;
  rom[15712] = 16'h10a1;
  rom[15713] = 16'h18c2;
  rom[15714] = 16'h18a2;
  rom[15715] = 16'h18c2;
  rom[15716] = 16'h18c2;
  rom[15717] = 16'h18c2;
  rom[15718] = 16'h18a2;
  rom[15719] = 16'h18c2;
  rom[15720] = 16'h10a1;
  rom[15721] = 16'h18c2;
  rom[15722] = 16'h0880;
  rom[15723] = 16'h20c3;
  rom[15724] = 16'h10c2;
  rom[15725] = 16'h6b4d;
  rom[15726] = 16'hef7d;
  rom[15727] = 16'hffff;
  rom[15728] = 16'hffdf;
  rom[15729] = 16'hffff;
  rom[15730] = 16'hffff;
  rom[15731] = 16'hffff;
  rom[15732] = 16'hffff;
  rom[15733] = 16'hffff;
  rom[15734] = 16'hffff;
  rom[15735] = 16'hffff;
  rom[15736] = 16'hffff;
  rom[15737] = 16'hffff;
  rom[15738] = 16'hffff;
  rom[15739] = 16'hffff;
  rom[15740] = 16'hffff;
  rom[15741] = 16'hb4d2;
  rom[15742] = 16'hbc6b;
  rom[15743] = 16'hed6a;
  rom[15744] = 16'hf549;
  rom[15745] = 16'hfd68;
  rom[15746] = 16'hfd47;
  rom[15747] = 16'hfd48;
  rom[15748] = 16'hfd28;
  rom[15749] = 16'hf529;
  rom[15750] = 16'hf529;
  rom[15751] = 16'hf528;
  rom[15752] = 16'he52b;
  rom[15753] = 16'habea;
  rom[15754] = 16'hd5d6;
  rom[15755] = 16'hffdf;
  rom[15756] = 16'hffff;
  rom[15757] = 16'hffff;
  rom[15758] = 16'hffff;
  rom[15759] = 16'hffff;
  rom[15760] = 16'hffff;
  rom[15761] = 16'hffff;
  rom[15762] = 16'hffff;
  rom[15763] = 16'hffff;
  rom[15764] = 16'hffff;
  rom[15765] = 16'hffff;
  rom[15766] = 16'hffff;
  rom[15767] = 16'hffff;
  rom[15768] = 16'hffff;
  rom[15769] = 16'hffff;
  rom[15770] = 16'hffff;
  rom[15771] = 16'hffff;
  rom[15772] = 16'hffff;
  rom[15773] = 16'hffff;
  rom[15774] = 16'hffff;
  rom[15775] = 16'hffff;
  rom[15776] = 16'hffff;
  rom[15777] = 16'hffff;
  rom[15778] = 16'hffff;
  rom[15779] = 16'hffff;
  rom[15780] = 16'hffff;
  rom[15781] = 16'hffff;
  rom[15782] = 16'hffff;
  rom[15783] = 16'hffff;
  rom[15784] = 16'hffff;
  rom[15785] = 16'hffff;
  rom[15786] = 16'hffff;
  rom[15787] = 16'hffff;
  rom[15788] = 16'hffff;
  rom[15789] = 16'hffff;
  rom[15790] = 16'hffff;
  rom[15791] = 16'hffff;
  rom[15792] = 16'hffff;
  rom[15793] = 16'hffff;
  rom[15794] = 16'hffff;
  rom[15795] = 16'hffff;
  rom[15796] = 16'hffff;
  rom[15797] = 16'hffff;
  rom[15798] = 16'hffff;
  rom[15799] = 16'hffff;
  rom[15800] = 16'hffff;
  rom[15801] = 16'hffff;
  rom[15802] = 16'hffff;
  rom[15803] = 16'hffff;
  rom[15804] = 16'hffff;
  rom[15805] = 16'hffff;
  rom[15806] = 16'hffff;
  rom[15807] = 16'hffff;
  rom[15808] = 16'hffff;
  rom[15809] = 16'hffff;
  rom[15810] = 16'hffff;
  rom[15811] = 16'hffff;
  rom[15812] = 16'hffff;
  rom[15813] = 16'hffff;
  rom[15814] = 16'hffff;
  rom[15815] = 16'hffff;
  rom[15816] = 16'hffff;
  rom[15817] = 16'hffff;
  rom[15818] = 16'hffff;
  rom[15819] = 16'hffff;
  rom[15820] = 16'hffff;
  rom[15821] = 16'hffff;
  rom[15822] = 16'hffff;
  rom[15823] = 16'hffff;
  rom[15824] = 16'hffff;
  rom[15825] = 16'hffff;
  rom[15826] = 16'hffff;
  rom[15827] = 16'hffff;
  rom[15828] = 16'hffff;
  rom[15829] = 16'hef19;
  rom[15830] = 16'h7ba8;
  rom[15831] = 16'h7bc5;
  rom[15832] = 16'he6ae;
  rom[15833] = 16'heecb;
  rom[15834] = 16'hff6c;
  rom[15835] = 16'hf709;
  rom[15836] = 16'hff2a;
  rom[15837] = 16'hff29;
  rom[15838] = 16'hf6e8;
  rom[15839] = 16'hf729;
  rom[15840] = 16'hff29;
  rom[15841] = 16'hf708;
  rom[15842] = 16'hf709;
  rom[15843] = 16'hff49;
  rom[15844] = 16'hff4a;
  rom[15845] = 16'hff4b;
  rom[15846] = 16'heeac;
  rom[15847] = 16'h7b03;
  rom[15848] = 16'h9b44;
  rom[15849] = 16'he52a;
  rom[15850] = 16'hfdab;
  rom[15851] = 16'he569;
  rom[15852] = 16'h72a5;
  rom[15853] = 16'hce18;
  rom[15854] = 16'hffff;
  rom[15855] = 16'hffff;
  rom[15856] = 16'hffff;
  rom[15857] = 16'hffff;
  rom[15858] = 16'hffff;
  rom[15859] = 16'hffff;
  rom[15860] = 16'hffff;
  rom[15861] = 16'hffff;
  rom[15862] = 16'hffff;
  rom[15863] = 16'hffff;
  rom[15864] = 16'hffff;
  rom[15865] = 16'hffff;
  rom[15866] = 16'hffff;
  rom[15867] = 16'hf77d;
  rom[15868] = 16'h6b4d;
  rom[15869] = 16'h18a2;
  rom[15870] = 16'h18a2;
  rom[15871] = 16'h10a1;
  rom[15872] = 16'h20e3;
  rom[15873] = 16'h10a1;
  rom[15874] = 16'h20e3;
  rom[15875] = 16'h18a2;
  rom[15876] = 16'h18c2;
  rom[15877] = 16'h18c2;
  rom[15878] = 16'h18a2;
  rom[15879] = 16'h18c2;
  rom[15880] = 16'h18a2;
  rom[15881] = 16'h18e3;
  rom[15882] = 16'h18c2;
  rom[15883] = 16'h18c3;
  rom[15884] = 16'h18a2;
  rom[15885] = 16'h18a2;
  rom[15886] = 16'h10a2;
  rom[15887] = 16'h18a1;
  rom[15888] = 16'h18a2;
  rom[15889] = 16'h6b4d;
  rom[15890] = 16'hffbf;
  rom[15891] = 16'hffff;
  rom[15892] = 16'hffff;
  rom[15893] = 16'hffff;
  rom[15894] = 16'hffff;
  rom[15895] = 16'hffff;
  rom[15896] = 16'hffff;
  rom[15897] = 16'hffff;
  rom[15898] = 16'hffff;
  rom[15899] = 16'hffff;
  rom[15900] = 16'hffff;
  rom[15901] = 16'hffff;
  rom[15902] = 16'hffff;
  rom[15903] = 16'hffff;
  rom[15904] = 16'hce39;
  rom[15905] = 16'h1082;
  rom[15906] = 16'h18c2;
  rom[15907] = 16'h18e3;
  rom[15908] = 16'h10a2;
  rom[15909] = 16'h18c2;
  rom[15910] = 16'h10a2;
  rom[15911] = 16'h18c2;
  rom[15912] = 16'h18c2;
  rom[15913] = 16'h10c2;
  rom[15914] = 16'h18c2;
  rom[15915] = 16'h18c2;
  rom[15916] = 16'h18c3;
  rom[15917] = 16'h18a2;
  rom[15918] = 16'h18a2;
  rom[15919] = 16'h20e3;
  rom[15920] = 16'h20c3;
  rom[15921] = 16'h1081;
  rom[15922] = 16'h18a2;
  rom[15923] = 16'h18c2;
  rom[15924] = 16'h18a2;
  rom[15925] = 16'h39a7;
  rom[15926] = 16'hc5d7;
  rom[15927] = 16'hffff;
  rom[15928] = 16'hffff;
  rom[15929] = 16'hffff;
  rom[15930] = 16'hffff;
  rom[15931] = 16'hffff;
  rom[15932] = 16'hffff;
  rom[15933] = 16'hffff;
  rom[15934] = 16'hffff;
  rom[15935] = 16'hffff;
  rom[15936] = 16'hffff;
  rom[15937] = 16'hffff;
  rom[15938] = 16'hffff;
  rom[15939] = 16'hffff;
  rom[15940] = 16'hffff;
  rom[15941] = 16'h9c0e;
  rom[15942] = 16'hc48b;
  rom[15943] = 16'hf54a;
  rom[15944] = 16'hfd49;
  rom[15945] = 16'hf547;
  rom[15946] = 16'hfd68;
  rom[15947] = 16'hfd47;
  rom[15948] = 16'hfd69;
  rom[15949] = 16'hf528;
  rom[15950] = 16'hfd69;
  rom[15951] = 16'hf508;
  rom[15952] = 16'hed4c;
  rom[15953] = 16'h9bca;
  rom[15954] = 16'hde37;
  rom[15955] = 16'hffff;
  rom[15956] = 16'hffff;
  rom[15957] = 16'hffff;
  rom[15958] = 16'hffff;
  rom[15959] = 16'hffff;
  rom[15960] = 16'hffff;
  rom[15961] = 16'hffff;
  rom[15962] = 16'hffff;
  rom[15963] = 16'hffff;
  rom[15964] = 16'hffff;
  rom[15965] = 16'hffff;
  rom[15966] = 16'hffff;
  rom[15967] = 16'hffff;
  rom[15968] = 16'hffff;
  rom[15969] = 16'hffff;
  rom[15970] = 16'hffff;
  rom[15971] = 16'hffff;
  rom[15972] = 16'hffff;
  rom[15973] = 16'hffff;
  rom[15974] = 16'hffff;
  rom[15975] = 16'hffff;
  rom[15976] = 16'hffff;
  rom[15977] = 16'hffff;
  rom[15978] = 16'hffff;
  rom[15979] = 16'hffff;
  rom[15980] = 16'hffff;
  rom[15981] = 16'hffff;
  rom[15982] = 16'hffff;
  rom[15983] = 16'hffff;
  rom[15984] = 16'hffff;
  rom[15985] = 16'hffff;
  rom[15986] = 16'hffff;
  rom[15987] = 16'hffff;
  rom[15988] = 16'hffff;
  rom[15989] = 16'hffff;
  rom[15990] = 16'hffff;
  rom[15991] = 16'hffff;
  rom[15992] = 16'hffff;
  rom[15993] = 16'hffff;
  rom[15994] = 16'hffff;
  rom[15995] = 16'hffff;
  rom[15996] = 16'hffff;
  rom[15997] = 16'hffff;
  rom[15998] = 16'hffff;
  rom[15999] = 16'hffff;
  rom[16000] = 16'hffff;
  rom[16001] = 16'hffff;
  rom[16002] = 16'hffff;
  rom[16003] = 16'hffff;
  rom[16004] = 16'hffff;
  rom[16005] = 16'hffff;
  rom[16006] = 16'hffff;
  rom[16007] = 16'hffff;
  rom[16008] = 16'hffff;
  rom[16009] = 16'hffff;
  rom[16010] = 16'hffff;
  rom[16011] = 16'hffff;
  rom[16012] = 16'hffff;
  rom[16013] = 16'hffff;
  rom[16014] = 16'hffff;
  rom[16015] = 16'hffff;
  rom[16016] = 16'hffff;
  rom[16017] = 16'hffff;
  rom[16018] = 16'hffff;
  rom[16019] = 16'hffff;
  rom[16020] = 16'hffff;
  rom[16021] = 16'hffff;
  rom[16022] = 16'hffff;
  rom[16023] = 16'hffff;
  rom[16024] = 16'hffff;
  rom[16025] = 16'hffff;
  rom[16026] = 16'hffdf;
  rom[16027] = 16'hffff;
  rom[16028] = 16'hf77b;
  rom[16029] = 16'h9cce;
  rom[16030] = 16'h7ba6;
  rom[16031] = 16'hde6d;
  rom[16032] = 16'hef0d;
  rom[16033] = 16'hf70b;
  rom[16034] = 16'hef09;
  rom[16035] = 16'hff29;
  rom[16036] = 16'hf728;
  rom[16037] = 16'hff29;
  rom[16038] = 16'hf708;
  rom[16039] = 16'hff29;
  rom[16040] = 16'hf708;
  rom[16041] = 16'hf729;
  rom[16042] = 16'hff29;
  rom[16043] = 16'hff29;
  rom[16044] = 16'hf709;
  rom[16045] = 16'hff29;
  rom[16046] = 16'hf6ec;
  rom[16047] = 16'hac87;
  rom[16048] = 16'h7281;
  rom[16049] = 16'he54b;
  rom[16050] = 16'hed27;
  rom[16051] = 16'hed8a;
  rom[16052] = 16'h9368;
  rom[16053] = 16'hbd75;
  rom[16054] = 16'hffdf;
  rom[16055] = 16'hffff;
  rom[16056] = 16'hffff;
  rom[16057] = 16'hffff;
  rom[16058] = 16'hffff;
  rom[16059] = 16'hffff;
  rom[16060] = 16'hffff;
  rom[16061] = 16'hffff;
  rom[16062] = 16'hffff;
  rom[16063] = 16'hffff;
  rom[16064] = 16'hffff;
  rom[16065] = 16'hffff;
  rom[16066] = 16'hffff;
  rom[16067] = 16'hd659;
  rom[16068] = 16'h31a5;
  rom[16069] = 16'h18e2;
  rom[16070] = 16'h1081;
  rom[16071] = 16'h20c3;
  rom[16072] = 16'h1081;
  rom[16073] = 16'h18c3;
  rom[16074] = 16'h18c2;
  rom[16075] = 16'h18c2;
  rom[16076] = 16'h10a1;
  rom[16077] = 16'h18c2;
  rom[16078] = 16'h18a2;
  rom[16079] = 16'h18c2;
  rom[16080] = 16'h10c2;
  rom[16081] = 16'h10a2;
  rom[16082] = 16'h10a2;
  rom[16083] = 16'h18c2;
  rom[16084] = 16'h18c2;
  rom[16085] = 16'h10a2;
  rom[16086] = 16'h10a2;
  rom[16087] = 16'h18c2;
  rom[16088] = 16'h1081;
  rom[16089] = 16'h3185;
  rom[16090] = 16'hd6ba;
  rom[16091] = 16'hffff;
  rom[16092] = 16'hffff;
  rom[16093] = 16'hffff;
  rom[16094] = 16'hffff;
  rom[16095] = 16'hffff;
  rom[16096] = 16'hffff;
  rom[16097] = 16'hffff;
  rom[16098] = 16'hffff;
  rom[16099] = 16'hffff;
  rom[16100] = 16'hffff;
  rom[16101] = 16'hffff;
  rom[16102] = 16'hffff;
  rom[16103] = 16'hffdf;
  rom[16104] = 16'h6b6d;
  rom[16105] = 16'h2103;
  rom[16106] = 16'h1081;
  rom[16107] = 16'h2103;
  rom[16108] = 16'h10a1;
  rom[16109] = 16'h10a1;
  rom[16110] = 16'h18c2;
  rom[16111] = 16'h1882;
  rom[16112] = 16'h18c2;
  rom[16113] = 16'h18c2;
  rom[16114] = 16'h1081;
  rom[16115] = 16'h18c2;
  rom[16116] = 16'h10a2;
  rom[16117] = 16'h20c3;
  rom[16118] = 16'h18c2;
  rom[16119] = 16'h18a2;
  rom[16120] = 16'h18c2;
  rom[16121] = 16'h18c2;
  rom[16122] = 16'h18a2;
  rom[16123] = 16'h18a2;
  rom[16124] = 16'h18c2;
  rom[16125] = 16'h18c2;
  rom[16126] = 16'h7bef;
  rom[16127] = 16'hf79e;
  rom[16128] = 16'hffdf;
  rom[16129] = 16'hffff;
  rom[16130] = 16'hffff;
  rom[16131] = 16'hffff;
  rom[16132] = 16'hffff;
  rom[16133] = 16'hffff;
  rom[16134] = 16'hffff;
  rom[16135] = 16'hffff;
  rom[16136] = 16'hffff;
  rom[16137] = 16'hffff;
  rom[16138] = 16'hffff;
  rom[16139] = 16'hffff;
  rom[16140] = 16'hffbe;
  rom[16141] = 16'h8329;
  rom[16142] = 16'hccab;
  rom[16143] = 16'hf54a;
  rom[16144] = 16'hf527;
  rom[16145] = 16'hfd68;
  rom[16146] = 16'hfd68;
  rom[16147] = 16'hfd67;
  rom[16148] = 16'hf548;
  rom[16149] = 16'hfd28;
  rom[16150] = 16'hfd28;
  rom[16151] = 16'hfd08;
  rom[16152] = 16'he50b;
  rom[16153] = 16'ha3ca;
  rom[16154] = 16'hce16;
  rom[16155] = 16'hffff;
  rom[16156] = 16'hffdf;
  rom[16157] = 16'hffff;
  rom[16158] = 16'hffff;
  rom[16159] = 16'hffff;
  rom[16160] = 16'hffff;
  rom[16161] = 16'hffff;
  rom[16162] = 16'hffff;
  rom[16163] = 16'hffff;
  rom[16164] = 16'hffff;
  rom[16165] = 16'hffff;
  rom[16166] = 16'hffff;
  rom[16167] = 16'hffff;
  rom[16168] = 16'hffff;
  rom[16169] = 16'hffff;
  rom[16170] = 16'hffff;
  rom[16171] = 16'hffff;
  rom[16172] = 16'hffff;
  rom[16173] = 16'hffff;
  rom[16174] = 16'hffff;
  rom[16175] = 16'hffff;
  rom[16176] = 16'hffff;
  rom[16177] = 16'hffff;
  rom[16178] = 16'hffff;
  rom[16179] = 16'hffff;
  rom[16180] = 16'hffff;
  rom[16181] = 16'hffff;
  rom[16182] = 16'hffff;
  rom[16183] = 16'hffff;
  rom[16184] = 16'hffff;
  rom[16185] = 16'hffff;
  rom[16186] = 16'hffff;
  rom[16187] = 16'hffff;
  rom[16188] = 16'hffff;
  rom[16189] = 16'hffff;
  rom[16190] = 16'hffff;
  rom[16191] = 16'hffff;
  rom[16192] = 16'hffff;
  rom[16193] = 16'hffff;
  rom[16194] = 16'hffff;
  rom[16195] = 16'hffff;
  rom[16196] = 16'hffff;
  rom[16197] = 16'hffff;
  rom[16198] = 16'hffff;
  rom[16199] = 16'hffff;
  rom[16200] = 16'hffff;
  rom[16201] = 16'hffff;
  rom[16202] = 16'hffff;
  rom[16203] = 16'hffff;
  rom[16204] = 16'hffff;
  rom[16205] = 16'hffff;
  rom[16206] = 16'hffff;
  rom[16207] = 16'hffff;
  rom[16208] = 16'hffff;
  rom[16209] = 16'hffff;
  rom[16210] = 16'hffff;
  rom[16211] = 16'hffff;
  rom[16212] = 16'hffff;
  rom[16213] = 16'hffff;
  rom[16214] = 16'hffff;
  rom[16215] = 16'hffff;
  rom[16216] = 16'hffff;
  rom[16217] = 16'hffff;
  rom[16218] = 16'hffff;
  rom[16219] = 16'hffff;
  rom[16220] = 16'hffff;
  rom[16221] = 16'hffff;
  rom[16222] = 16'hffff;
  rom[16223] = 16'hffff;
  rom[16224] = 16'hffff;
  rom[16225] = 16'hffff;
  rom[16226] = 16'hffbf;
  rom[16227] = 16'hffde;
  rom[16228] = 16'hdeb8;
  rom[16229] = 16'h4a41;
  rom[16230] = 16'hc5ac;
  rom[16231] = 16'hff6f;
  rom[16232] = 16'hff4d;
  rom[16233] = 16'hff4b;
  rom[16234] = 16'hf6e8;
  rom[16235] = 16'hff29;
  rom[16236] = 16'hff29;
  rom[16237] = 16'hff29;
  rom[16238] = 16'hf6e9;
  rom[16239] = 16'hff49;
  rom[16240] = 16'hff2a;
  rom[16241] = 16'hf728;
  rom[16242] = 16'hff4a;
  rom[16243] = 16'hff29;
  rom[16244] = 16'hff4a;
  rom[16245] = 16'hff49;
  rom[16246] = 16'hff0c;
  rom[16247] = 16'hc569;
  rom[16248] = 16'h6a02;
  rom[16249] = 16'hd4e8;
  rom[16250] = 16'hfdca;
  rom[16251] = 16'hed49;
  rom[16252] = 16'hb42a;
  rom[16253] = 16'h8bed;
  rom[16254] = 16'hffff;
  rom[16255] = 16'hffff;
  rom[16256] = 16'hffff;
  rom[16257] = 16'hffff;
  rom[16258] = 16'hffff;
  rom[16259] = 16'hffff;
  rom[16260] = 16'hffff;
  rom[16261] = 16'hffff;
  rom[16262] = 16'hffff;
  rom[16263] = 16'hffff;
  rom[16264] = 16'hffff;
  rom[16265] = 16'hffff;
  rom[16266] = 16'hffff;
  rom[16267] = 16'hb575;
  rom[16268] = 16'h20e3;
  rom[16269] = 16'h18a2;
  rom[16270] = 16'h2103;
  rom[16271] = 16'h18a2;
  rom[16272] = 16'h10a2;
  rom[16273] = 16'h10a1;
  rom[16274] = 16'h18e3;
  rom[16275] = 16'h10a1;
  rom[16276] = 16'h18e2;
  rom[16277] = 16'h18c2;
  rom[16278] = 16'h20e3;
  rom[16279] = 16'h18c2;
  rom[16280] = 16'h5acb;
  rom[16281] = 16'had55;
  rom[16282] = 16'hb555;
  rom[16283] = 16'h5acb;
  rom[16284] = 16'h20e3;
  rom[16285] = 16'h18c2;
  rom[16286] = 16'h18c2;
  rom[16287] = 16'h18c2;
  rom[16288] = 16'h2103;
  rom[16289] = 16'h10a1;
  rom[16290] = 16'hbdd6;
  rom[16291] = 16'hffff;
  rom[16292] = 16'hffff;
  rom[16293] = 16'hffff;
  rom[16294] = 16'hffff;
  rom[16295] = 16'hffff;
  rom[16296] = 16'hffff;
  rom[16297] = 16'hffff;
  rom[16298] = 16'hffff;
  rom[16299] = 16'hffff;
  rom[16300] = 16'hffff;
  rom[16301] = 16'hffff;
  rom[16302] = 16'hffff;
  rom[16303] = 16'he6fb;
  rom[16304] = 16'h4a28;
  rom[16305] = 16'h18c3;
  rom[16306] = 16'h10a2;
  rom[16307] = 16'h1081;
  rom[16308] = 16'h20e3;
  rom[16309] = 16'h10a2;
  rom[16310] = 16'h4a08;
  rom[16311] = 16'h8c51;
  rom[16312] = 16'had14;
  rom[16313] = 16'h6b8d;
  rom[16314] = 16'h4208;
  rom[16315] = 16'h0861;
  rom[16316] = 16'h2124;
  rom[16317] = 16'h1061;
  rom[16318] = 16'h20c3;
  rom[16319] = 16'h18a2;
  rom[16320] = 16'h18a2;
  rom[16321] = 16'h18a2;
  rom[16322] = 16'h18a2;
  rom[16323] = 16'h18c2;
  rom[16324] = 16'h10c2;
  rom[16325] = 16'h18e3;
  rom[16326] = 16'h31a6;
  rom[16327] = 16'he6fb;
  rom[16328] = 16'hffff;
  rom[16329] = 16'hffff;
  rom[16330] = 16'hffff;
  rom[16331] = 16'hffff;
  rom[16332] = 16'hffff;
  rom[16333] = 16'hffff;
  rom[16334] = 16'hffff;
  rom[16335] = 16'hffff;
  rom[16336] = 16'hffff;
  rom[16337] = 16'hffff;
  rom[16338] = 16'hffff;
  rom[16339] = 16'hffff;
  rom[16340] = 16'hf75c;
  rom[16341] = 16'h72c7;
  rom[16342] = 16'hd4ec;
  rom[16343] = 16'hf529;
  rom[16344] = 16'hfd49;
  rom[16345] = 16'hfd28;
  rom[16346] = 16'hfd68;
  rom[16347] = 16'hf527;
  rom[16348] = 16'hfd48;
  rom[16349] = 16'hf528;
  rom[16350] = 16'hfd28;
  rom[16351] = 16'hfd28;
  rom[16352] = 16'hed4c;
  rom[16353] = 16'ha3ca;
  rom[16354] = 16'hde18;
  rom[16355] = 16'hffff;
  rom[16356] = 16'hffff;
  rom[16357] = 16'hffff;
  rom[16358] = 16'hffff;
  rom[16359] = 16'hffff;
  rom[16360] = 16'hffff;
  rom[16361] = 16'hffff;
  rom[16362] = 16'hffff;
  rom[16363] = 16'hffff;
  rom[16364] = 16'hffff;
  rom[16365] = 16'hffff;
  rom[16366] = 16'hffff;
  rom[16367] = 16'hffff;
  rom[16368] = 16'hffff;
  rom[16369] = 16'hffff;
  rom[16370] = 16'hffff;
  rom[16371] = 16'hffff;
  rom[16372] = 16'hffff;
  rom[16373] = 16'hffff;
  rom[16374] = 16'hffff;
  rom[16375] = 16'hffff;
  rom[16376] = 16'hffff;
  rom[16377] = 16'hffff;
  rom[16378] = 16'hffff;
  rom[16379] = 16'hffff;
  rom[16380] = 16'hffff;
  rom[16381] = 16'hffff;
  rom[16382] = 16'hffff;
  rom[16383] = 16'hffff;
  rom[16384] = 16'hffff;
  rom[16385] = 16'hffff;
  rom[16386] = 16'hffff;
  rom[16387] = 16'hffff;
  rom[16388] = 16'hffff;
  rom[16389] = 16'hffff;
  rom[16390] = 16'hffff;
  rom[16391] = 16'hffff;
  rom[16392] = 16'hffff;
  rom[16393] = 16'hffff;
  rom[16394] = 16'hffff;
  rom[16395] = 16'hffff;
  rom[16396] = 16'hffff;
  rom[16397] = 16'hffff;
  rom[16398] = 16'hffff;
  rom[16399] = 16'hffff;
  rom[16400] = 16'hffff;
  rom[16401] = 16'hffff;
  rom[16402] = 16'hffff;
  rom[16403] = 16'hffff;
  rom[16404] = 16'hffff;
  rom[16405] = 16'hffff;
  rom[16406] = 16'hffff;
  rom[16407] = 16'hffff;
  rom[16408] = 16'hffff;
  rom[16409] = 16'hffff;
  rom[16410] = 16'hffff;
  rom[16411] = 16'hffff;
  rom[16412] = 16'hffff;
  rom[16413] = 16'hffff;
  rom[16414] = 16'hffff;
  rom[16415] = 16'hffff;
  rom[16416] = 16'hffff;
  rom[16417] = 16'hffff;
  rom[16418] = 16'hffff;
  rom[16419] = 16'hffff;
  rom[16420] = 16'hffff;
  rom[16421] = 16'hffff;
  rom[16422] = 16'hffff;
  rom[16423] = 16'hffff;
  rom[16424] = 16'hffff;
  rom[16425] = 16'hffdf;
  rom[16426] = 16'hffff;
  rom[16427] = 16'hf75c;
  rom[16428] = 16'h83aa;
  rom[16429] = 16'h83a5;
  rom[16430] = 16'he6cc;
  rom[16431] = 16'hf72c;
  rom[16432] = 16'heee9;
  rom[16433] = 16'hff2a;
  rom[16434] = 16'hf708;
  rom[16435] = 16'hff28;
  rom[16436] = 16'hf728;
  rom[16437] = 16'hff29;
  rom[16438] = 16'hf728;
  rom[16439] = 16'hff28;
  rom[16440] = 16'hff28;
  rom[16441] = 16'hff29;
  rom[16442] = 16'hf708;
  rom[16443] = 16'hff29;
  rom[16444] = 16'hf708;
  rom[16445] = 16'hff49;
  rom[16446] = 16'hf70a;
  rom[16447] = 16'hc569;
  rom[16448] = 16'h69e1;
  rom[16449] = 16'hdce9;
  rom[16450] = 16'hf568;
  rom[16451] = 16'hf549;
  rom[16452] = 16'hc46a;
  rom[16453] = 16'h830a;
  rom[16454] = 16'hff9e;
  rom[16455] = 16'hffff;
  rom[16456] = 16'hffff;
  rom[16457] = 16'hffff;
  rom[16458] = 16'hffff;
  rom[16459] = 16'hffff;
  rom[16460] = 16'hffff;
  rom[16461] = 16'hffff;
  rom[16462] = 16'hffff;
  rom[16463] = 16'hffff;
  rom[16464] = 16'hffff;
  rom[16465] = 16'hffff;
  rom[16466] = 16'hffbe;
  rom[16467] = 16'h7bef;
  rom[16468] = 16'h18c2;
  rom[16469] = 16'h18a2;
  rom[16470] = 16'h10a2;
  rom[16471] = 16'h18c3;
  rom[16472] = 16'h10a1;
  rom[16473] = 16'h18c2;
  rom[16474] = 16'h10a2;
  rom[16475] = 16'h18c2;
  rom[16476] = 16'h18c2;
  rom[16477] = 16'h18a2;
  rom[16478] = 16'h2964;
  rom[16479] = 16'hb596;
  rom[16480] = 16'hf79e;
  rom[16481] = 16'hffff;
  rom[16482] = 16'hffdf;
  rom[16483] = 16'hffdf;
  rom[16484] = 16'hc618;
  rom[16485] = 16'h4a69;
  rom[16486] = 16'h10a2;
  rom[16487] = 16'h10a2;
  rom[16488] = 16'h18c3;
  rom[16489] = 16'h18a2;
  rom[16490] = 16'h8410;
  rom[16491] = 16'hffff;
  rom[16492] = 16'hffff;
  rom[16493] = 16'hffff;
  rom[16494] = 16'hffff;
  rom[16495] = 16'hffff;
  rom[16496] = 16'hffff;
  rom[16497] = 16'hffff;
  rom[16498] = 16'hffff;
  rom[16499] = 16'hffff;
  rom[16500] = 16'hffff;
  rom[16501] = 16'hffff;
  rom[16502] = 16'hffff;
  rom[16503] = 16'hdebb;
  rom[16504] = 16'h2965;
  rom[16505] = 16'h10a2;
  rom[16506] = 16'h18c2;
  rom[16507] = 16'h1082;
  rom[16508] = 16'h2944;
  rom[16509] = 16'h8c51;
  rom[16510] = 16'hef5d;
  rom[16511] = 16'hffdf;
  rom[16512] = 16'hffff;
  rom[16513] = 16'hffff;
  rom[16514] = 16'hd69a;
  rom[16515] = 16'h83ef;
  rom[16516] = 16'h10c2;
  rom[16517] = 16'h20e3;
  rom[16518] = 16'h18a2;
  rom[16519] = 16'h18c2;
  rom[16520] = 16'h18a2;
  rom[16521] = 16'h18c3;
  rom[16522] = 16'h18a2;
  rom[16523] = 16'h18c2;
  rom[16524] = 16'h10a2;
  rom[16525] = 16'h10a2;
  rom[16526] = 16'h20e3;
  rom[16527] = 16'hd679;
  rom[16528] = 16'hffff;
  rom[16529] = 16'hffff;
  rom[16530] = 16'hffff;
  rom[16531] = 16'hffff;
  rom[16532] = 16'hffff;
  rom[16533] = 16'hffff;
  rom[16534] = 16'hffff;
  rom[16535] = 16'hffff;
  rom[16536] = 16'hffff;
  rom[16537] = 16'hffff;
  rom[16538] = 16'hfffe;
  rom[16539] = 16'hffff;
  rom[16540] = 16'hd637;
  rom[16541] = 16'h8b48;
  rom[16542] = 16'hdd0a;
  rom[16543] = 16'hf549;
  rom[16544] = 16'hfd28;
  rom[16545] = 16'hfd29;
  rom[16546] = 16'hf528;
  rom[16547] = 16'hfd47;
  rom[16548] = 16'hf548;
  rom[16549] = 16'hfd28;
  rom[16550] = 16'hf4e6;
  rom[16551] = 16'hfd28;
  rom[16552] = 16'he52b;
  rom[16553] = 16'h9369;
  rom[16554] = 16'hce16;
  rom[16555] = 16'hffff;
  rom[16556] = 16'hffff;
  rom[16557] = 16'hffff;
  rom[16558] = 16'hffff;
  rom[16559] = 16'hffff;
  rom[16560] = 16'hffff;
  rom[16561] = 16'hffff;
  rom[16562] = 16'hffff;
  rom[16563] = 16'hffff;
  rom[16564] = 16'hffff;
  rom[16565] = 16'hffff;
  rom[16566] = 16'hffff;
  rom[16567] = 16'hffff;
  rom[16568] = 16'hffff;
  rom[16569] = 16'hffff;
  rom[16570] = 16'hffff;
  rom[16571] = 16'hffff;
  rom[16572] = 16'hffff;
  rom[16573] = 16'hffff;
  rom[16574] = 16'hffff;
  rom[16575] = 16'hffff;
  rom[16576] = 16'hffff;
  rom[16577] = 16'hffff;
  rom[16578] = 16'hffff;
  rom[16579] = 16'hffff;
  rom[16580] = 16'hffff;
  rom[16581] = 16'hffff;
  rom[16582] = 16'hffff;
  rom[16583] = 16'hffff;
  rom[16584] = 16'hffff;
  rom[16585] = 16'hffff;
  rom[16586] = 16'hffff;
  rom[16587] = 16'hffff;
  rom[16588] = 16'hffff;
  rom[16589] = 16'hffff;
  rom[16590] = 16'hffff;
  rom[16591] = 16'hffff;
  rom[16592] = 16'hffff;
  rom[16593] = 16'hffff;
  rom[16594] = 16'hffff;
  rom[16595] = 16'hffff;
  rom[16596] = 16'hffff;
  rom[16597] = 16'hffff;
  rom[16598] = 16'hffff;
  rom[16599] = 16'hffff;
  rom[16600] = 16'hffff;
  rom[16601] = 16'hffff;
  rom[16602] = 16'hffff;
  rom[16603] = 16'hffff;
  rom[16604] = 16'hffff;
  rom[16605] = 16'hffff;
  rom[16606] = 16'hffff;
  rom[16607] = 16'hffff;
  rom[16608] = 16'hffff;
  rom[16609] = 16'hffff;
  rom[16610] = 16'hffff;
  rom[16611] = 16'hffff;
  rom[16612] = 16'hffff;
  rom[16613] = 16'hffff;
  rom[16614] = 16'hffff;
  rom[16615] = 16'hffff;
  rom[16616] = 16'hffff;
  rom[16617] = 16'hffff;
  rom[16618] = 16'hffff;
  rom[16619] = 16'hffff;
  rom[16620] = 16'hffff;
  rom[16621] = 16'hffff;
  rom[16622] = 16'hffff;
  rom[16623] = 16'hffff;
  rom[16624] = 16'hffff;
  rom[16625] = 16'hffdf;
  rom[16626] = 16'hffdf;
  rom[16627] = 16'he6b9;
  rom[16628] = 16'h6ae6;
  rom[16629] = 16'hcdcc;
  rom[16630] = 16'hff4d;
  rom[16631] = 16'hf6e8;
  rom[16632] = 16'hff4a;
  rom[16633] = 16'hff2a;
  rom[16634] = 16'hff29;
  rom[16635] = 16'hf708;
  rom[16636] = 16'hff49;
  rom[16637] = 16'hf728;
  rom[16638] = 16'hff49;
  rom[16639] = 16'hf729;
  rom[16640] = 16'hff29;
  rom[16641] = 16'hff29;
  rom[16642] = 16'hff49;
  rom[16643] = 16'hff29;
  rom[16644] = 16'hf709;
  rom[16645] = 16'hf708;
  rom[16646] = 16'hff4c;
  rom[16647] = 16'hb4c5;
  rom[16648] = 16'h7a62;
  rom[16649] = 16'hdce8;
  rom[16650] = 16'hfd89;
  rom[16651] = 16'hf549;
  rom[16652] = 16'hdd0d;
  rom[16653] = 16'h8308;
  rom[16654] = 16'heedb;
  rom[16655] = 16'hffff;
  rom[16656] = 16'hffff;
  rom[16657] = 16'hffff;
  rom[16658] = 16'hffff;
  rom[16659] = 16'hffff;
  rom[16660] = 16'hffff;
  rom[16661] = 16'hffff;
  rom[16662] = 16'hffff;
  rom[16663] = 16'hffff;
  rom[16664] = 16'hffff;
  rom[16665] = 16'hffff;
  rom[16666] = 16'hf79e;
  rom[16667] = 16'h528a;
  rom[16668] = 16'h20e3;
  rom[16669] = 16'h20e3;
  rom[16670] = 16'h18a2;
  rom[16671] = 16'h18c3;
  rom[16672] = 16'h18a2;
  rom[16673] = 16'h10a1;
  rom[16674] = 16'h18c3;
  rom[16675] = 16'h1081;
  rom[16676] = 16'h2904;
  rom[16677] = 16'h20e3;
  rom[16678] = 16'hbdd6;
  rom[16679] = 16'hffff;
  rom[16680] = 16'hffff;
  rom[16681] = 16'hffdf;
  rom[16682] = 16'hffff;
  rom[16683] = 16'hef7d;
  rom[16684] = 16'hffff;
  rom[16685] = 16'hc5f7;
  rom[16686] = 16'h3185;
  rom[16687] = 16'h1081;
  rom[16688] = 16'h20e3;
  rom[16689] = 16'h18c2;
  rom[16690] = 16'h5aca;
  rom[16691] = 16'hffdf;
  rom[16692] = 16'hffff;
  rom[16693] = 16'hffff;
  rom[16694] = 16'hffff;
  rom[16695] = 16'hffff;
  rom[16696] = 16'hffff;
  rom[16697] = 16'hffff;
  rom[16698] = 16'hffff;
  rom[16699] = 16'hffff;
  rom[16700] = 16'hffff;
  rom[16701] = 16'hffff;
  rom[16702] = 16'hffff;
  rom[16703] = 16'hce79;
  rom[16704] = 16'h2945;
  rom[16705] = 16'h2104;
  rom[16706] = 16'h18e3;
  rom[16707] = 16'h18a2;
  rom[16708] = 16'h83cf;
  rom[16709] = 16'hf79e;
  rom[16710] = 16'hffff;
  rom[16711] = 16'hffff;
  rom[16712] = 16'hffff;
  rom[16713] = 16'hffff;
  rom[16714] = 16'hffff;
  rom[16715] = 16'hdefb;
  rom[16716] = 16'h5269;
  rom[16717] = 16'h1041;
  rom[16718] = 16'h20e3;
  rom[16719] = 16'h1082;
  rom[16720] = 16'h18c2;
  rom[16721] = 16'h1082;
  rom[16722] = 16'h18c2;
  rom[16723] = 16'h18c2;
  rom[16724] = 16'h18c3;
  rom[16725] = 16'h10a2;
  rom[16726] = 16'h18e3;
  rom[16727] = 16'hc638;
  rom[16728] = 16'hffdf;
  rom[16729] = 16'hffff;
  rom[16730] = 16'hffff;
  rom[16731] = 16'hffff;
  rom[16732] = 16'hffff;
  rom[16733] = 16'hffff;
  rom[16734] = 16'hffff;
  rom[16735] = 16'hffff;
  rom[16736] = 16'hffff;
  rom[16737] = 16'hffff;
  rom[16738] = 16'hffff;
  rom[16739] = 16'hfffe;
  rom[16740] = 16'hacf1;
  rom[16741] = 16'h9bc9;
  rom[16742] = 16'he56b;
  rom[16743] = 16'hf548;
  rom[16744] = 16'hfd49;
  rom[16745] = 16'hfd29;
  rom[16746] = 16'hfd29;
  rom[16747] = 16'hfd48;
  rom[16748] = 16'hfd49;
  rom[16749] = 16'hfd28;
  rom[16750] = 16'hfce6;
  rom[16751] = 16'hfd28;
  rom[16752] = 16'he52c;
  rom[16753] = 16'h8307;
  rom[16754] = 16'hd637;
  rom[16755] = 16'hffff;
  rom[16756] = 16'hffff;
  rom[16757] = 16'hffff;
  rom[16758] = 16'hffff;
  rom[16759] = 16'hffff;
  rom[16760] = 16'hffff;
  rom[16761] = 16'hffff;
  rom[16762] = 16'hffff;
  rom[16763] = 16'hffff;
  rom[16764] = 16'hffff;
  rom[16765] = 16'hffff;
  rom[16766] = 16'hffff;
  rom[16767] = 16'hffff;
  rom[16768] = 16'hffff;
  rom[16769] = 16'hffff;
  rom[16770] = 16'hffff;
  rom[16771] = 16'hffff;
  rom[16772] = 16'hffff;
  rom[16773] = 16'hffff;
  rom[16774] = 16'hffff;
  rom[16775] = 16'hffff;
  rom[16776] = 16'hffff;
  rom[16777] = 16'hffff;
  rom[16778] = 16'hffff;
  rom[16779] = 16'hffff;
  rom[16780] = 16'hffff;
  rom[16781] = 16'hffff;
  rom[16782] = 16'hffff;
  rom[16783] = 16'hffff;
  rom[16784] = 16'hffff;
  rom[16785] = 16'hffff;
  rom[16786] = 16'hffff;
  rom[16787] = 16'hffff;
  rom[16788] = 16'hffff;
  rom[16789] = 16'hffff;
  rom[16790] = 16'hffff;
  rom[16791] = 16'hffff;
  rom[16792] = 16'hffff;
  rom[16793] = 16'hffff;
  rom[16794] = 16'hffff;
  rom[16795] = 16'hffff;
  rom[16796] = 16'hffff;
  rom[16797] = 16'hffff;
  rom[16798] = 16'hffff;
  rom[16799] = 16'hffff;
  rom[16800] = 16'hffff;
  rom[16801] = 16'hffff;
  rom[16802] = 16'hffff;
  rom[16803] = 16'hffff;
  rom[16804] = 16'hffff;
  rom[16805] = 16'hffff;
  rom[16806] = 16'hffff;
  rom[16807] = 16'hffff;
  rom[16808] = 16'hffff;
  rom[16809] = 16'hffff;
  rom[16810] = 16'hffff;
  rom[16811] = 16'hffff;
  rom[16812] = 16'hffff;
  rom[16813] = 16'hffff;
  rom[16814] = 16'hffff;
  rom[16815] = 16'hffff;
  rom[16816] = 16'hffff;
  rom[16817] = 16'hffff;
  rom[16818] = 16'hffff;
  rom[16819] = 16'hffff;
  rom[16820] = 16'hffff;
  rom[16821] = 16'hffff;
  rom[16822] = 16'hffff;
  rom[16823] = 16'hffff;
  rom[16824] = 16'hffdf;
  rom[16825] = 16'hffff;
  rom[16826] = 16'hffbe;
  rom[16827] = 16'hbdb4;
  rom[16828] = 16'h6b24;
  rom[16829] = 16'heeee;
  rom[16830] = 16'hf70a;
  rom[16831] = 16'hff28;
  rom[16832] = 16'hf709;
  rom[16833] = 16'hff2a;
  rom[16834] = 16'hf708;
  rom[16835] = 16'hff48;
  rom[16836] = 16'hf708;
  rom[16837] = 16'hff28;
  rom[16838] = 16'hff28;
  rom[16839] = 16'hff29;
  rom[16840] = 16'hf708;
  rom[16841] = 16'hff28;
  rom[16842] = 16'hff09;
  rom[16843] = 16'hff29;
  rom[16844] = 16'hf729;
  rom[16845] = 16'hf749;
  rom[16846] = 16'hf70a;
  rom[16847] = 16'hac84;
  rom[16848] = 16'h7241;
  rom[16849] = 16'he529;
  rom[16850] = 16'hf567;
  rom[16851] = 16'hf54a;
  rom[16852] = 16'hdd2c;
  rom[16853] = 16'h9369;
  rom[16854] = 16'hd617;
  rom[16855] = 16'hffdf;
  rom[16856] = 16'hffff;
  rom[16857] = 16'hffff;
  rom[16858] = 16'hffff;
  rom[16859] = 16'hffff;
  rom[16860] = 16'hffff;
  rom[16861] = 16'hffff;
  rom[16862] = 16'hffff;
  rom[16863] = 16'hffff;
  rom[16864] = 16'hffff;
  rom[16865] = 16'hffff;
  rom[16866] = 16'hf77e;
  rom[16867] = 16'h4a49;
  rom[16868] = 16'h18a2;
  rom[16869] = 16'h18c3;
  rom[16870] = 16'h18a2;
  rom[16871] = 16'h18a2;
  rom[16872] = 16'h18c2;
  rom[16873] = 16'h18a2;
  rom[16874] = 16'h18a2;
  rom[16875] = 16'h18c2;
  rom[16876] = 16'h0861;
  rom[16877] = 16'h39c6;
  rom[16878] = 16'hdefa;
  rom[16879] = 16'hffff;
  rom[16880] = 16'hffff;
  rom[16881] = 16'hffff;
  rom[16882] = 16'hffff;
  rom[16883] = 16'hffff;
  rom[16884] = 16'hffff;
  rom[16885] = 16'hf79e;
  rom[16886] = 16'h630b;
  rom[16887] = 16'h18e3;
  rom[16888] = 16'h18a2;
  rom[16889] = 16'h18c2;
  rom[16890] = 16'h4a48;
  rom[16891] = 16'hffdf;
  rom[16892] = 16'hffff;
  rom[16893] = 16'hffff;
  rom[16894] = 16'hffff;
  rom[16895] = 16'hffff;
  rom[16896] = 16'hffff;
  rom[16897] = 16'hffff;
  rom[16898] = 16'hffff;
  rom[16899] = 16'hffff;
  rom[16900] = 16'hffff;
  rom[16901] = 16'hffff;
  rom[16902] = 16'hffff;
  rom[16903] = 16'hd679;
  rom[16904] = 16'h2124;
  rom[16905] = 16'h10a2;
  rom[16906] = 16'h10a2;
  rom[16907] = 16'h2924;
  rom[16908] = 16'ha534;
  rom[16909] = 16'hffff;
  rom[16910] = 16'hffff;
  rom[16911] = 16'hffff;
  rom[16912] = 16'hffff;
  rom[16913] = 16'hffff;
  rom[16914] = 16'hffdf;
  rom[16915] = 16'hffdf;
  rom[16916] = 16'h8430;
  rom[16917] = 16'h18a2;
  rom[16918] = 16'h18c2;
  rom[16919] = 16'h1061;
  rom[16920] = 16'h18c2;
  rom[16921] = 16'h18a2;
  rom[16922] = 16'h18c2;
  rom[16923] = 16'h18c2;
  rom[16924] = 16'h10a2;
  rom[16925] = 16'h18c2;
  rom[16926] = 16'h18e3;
  rom[16927] = 16'hce39;
  rom[16928] = 16'hffff;
  rom[16929] = 16'hffdf;
  rom[16930] = 16'hffff;
  rom[16931] = 16'hffff;
  rom[16932] = 16'hffff;
  rom[16933] = 16'hffff;
  rom[16934] = 16'hffff;
  rom[16935] = 16'hffff;
  rom[16936] = 16'hffff;
  rom[16937] = 16'hffff;
  rom[16938] = 16'hffff;
  rom[16939] = 16'hff9d;
  rom[16940] = 16'h83aa;
  rom[16941] = 16'hac29;
  rom[16942] = 16'he56a;
  rom[16943] = 16'hf568;
  rom[16944] = 16'hfd27;
  rom[16945] = 16'hfd49;
  rom[16946] = 16'hf508;
  rom[16947] = 16'hfd48;
  rom[16948] = 16'hf528;
  rom[16949] = 16'hfd28;
  rom[16950] = 16'hfcc6;
  rom[16951] = 16'hfd49;
  rom[16952] = 16'hdd2c;
  rom[16953] = 16'h7b07;
  rom[16954] = 16'hde98;
  rom[16955] = 16'hffff;
  rom[16956] = 16'hffff;
  rom[16957] = 16'hffff;
  rom[16958] = 16'hffff;
  rom[16959] = 16'hffff;
  rom[16960] = 16'hffff;
  rom[16961] = 16'hffff;
  rom[16962] = 16'hffff;
  rom[16963] = 16'hffff;
  rom[16964] = 16'hffff;
  rom[16965] = 16'hffff;
  rom[16966] = 16'hffff;
  rom[16967] = 16'hffff;
  rom[16968] = 16'hffff;
  rom[16969] = 16'hffff;
  rom[16970] = 16'hffff;
  rom[16971] = 16'hffff;
  rom[16972] = 16'hffff;
  rom[16973] = 16'hffff;
  rom[16974] = 16'hffff;
  rom[16975] = 16'hffff;
  rom[16976] = 16'hffff;
  rom[16977] = 16'hffff;
  rom[16978] = 16'hffff;
  rom[16979] = 16'hffff;
  rom[16980] = 16'hffff;
  rom[16981] = 16'hffff;
  rom[16982] = 16'hffff;
  rom[16983] = 16'hffff;
  rom[16984] = 16'hffff;
  rom[16985] = 16'hffff;
  rom[16986] = 16'hffff;
  rom[16987] = 16'hffff;
  rom[16988] = 16'hffff;
  rom[16989] = 16'hffff;
  rom[16990] = 16'hffff;
  rom[16991] = 16'hffff;
  rom[16992] = 16'hffff;
  rom[16993] = 16'hffff;
  rom[16994] = 16'hffff;
  rom[16995] = 16'hffff;
  rom[16996] = 16'hffff;
  rom[16997] = 16'hffff;
  rom[16998] = 16'hffff;
  rom[16999] = 16'hffff;
  rom[17000] = 16'hffff;
  rom[17001] = 16'hffff;
  rom[17002] = 16'hffff;
  rom[17003] = 16'hffff;
  rom[17004] = 16'hffff;
  rom[17005] = 16'hffff;
  rom[17006] = 16'hffff;
  rom[17007] = 16'hffff;
  rom[17008] = 16'hffff;
  rom[17009] = 16'hffff;
  rom[17010] = 16'hffff;
  rom[17011] = 16'hffff;
  rom[17012] = 16'hffff;
  rom[17013] = 16'hffff;
  rom[17014] = 16'hffff;
  rom[17015] = 16'hffff;
  rom[17016] = 16'hffff;
  rom[17017] = 16'hffff;
  rom[17018] = 16'hffff;
  rom[17019] = 16'hffff;
  rom[17020] = 16'hffff;
  rom[17021] = 16'hffff;
  rom[17022] = 16'hffff;
  rom[17023] = 16'hffff;
  rom[17024] = 16'hffff;
  rom[17025] = 16'hffff;
  rom[17026] = 16'hffff;
  rom[17027] = 16'h9cce;
  rom[17028] = 16'h9c68;
  rom[17029] = 16'hf74e;
  rom[17030] = 16'hff4a;
  rom[17031] = 16'hff29;
  rom[17032] = 16'hff2a;
  rom[17033] = 16'hf6e9;
  rom[17034] = 16'hff49;
  rom[17035] = 16'hff28;
  rom[17036] = 16'hff29;
  rom[17037] = 16'hff28;
  rom[17038] = 16'hff29;
  rom[17039] = 16'hff28;
  rom[17040] = 16'hff29;
  rom[17041] = 16'hff28;
  rom[17042] = 16'hff29;
  rom[17043] = 16'hff29;
  rom[17044] = 16'hff2a;
  rom[17045] = 16'hf72a;
  rom[17046] = 16'hf6ea;
  rom[17047] = 16'ha422;
  rom[17048] = 16'h7a62;
  rom[17049] = 16'he54a;
  rom[17050] = 16'hf548;
  rom[17051] = 16'hf54a;
  rom[17052] = 16'hed6c;
  rom[17053] = 16'ha3e9;
  rom[17054] = 16'hacb0;
  rom[17055] = 16'hffdf;
  rom[17056] = 16'hffdf;
  rom[17057] = 16'hffff;
  rom[17058] = 16'hffff;
  rom[17059] = 16'hffff;
  rom[17060] = 16'hffff;
  rom[17061] = 16'hffff;
  rom[17062] = 16'hffff;
  rom[17063] = 16'hffff;
  rom[17064] = 16'hffff;
  rom[17065] = 16'hffdf;
  rom[17066] = 16'hffdf;
  rom[17067] = 16'h52aa;
  rom[17068] = 16'h18a2;
  rom[17069] = 16'h18a2;
  rom[17070] = 16'h20c3;
  rom[17071] = 16'h20c3;
  rom[17072] = 16'h18a2;
  rom[17073] = 16'h18a2;
  rom[17074] = 16'h20c3;
  rom[17075] = 16'h18a2;
  rom[17076] = 16'h2904;
  rom[17077] = 16'h41e7;
  rom[17078] = 16'hef5d;
  rom[17079] = 16'hffff;
  rom[17080] = 16'hffff;
  rom[17081] = 16'hffff;
  rom[17082] = 16'hffff;
  rom[17083] = 16'hffff;
  rom[17084] = 16'hffff;
  rom[17085] = 16'hffff;
  rom[17086] = 16'h83ef;
  rom[17087] = 16'h18a2;
  rom[17088] = 16'h18e3;
  rom[17089] = 16'h10a1;
  rom[17090] = 16'h630c;
  rom[17091] = 16'hffbf;
  rom[17092] = 16'hffff;
  rom[17093] = 16'hffff;
  rom[17094] = 16'hffff;
  rom[17095] = 16'hffff;
  rom[17096] = 16'hffff;
  rom[17097] = 16'hffff;
  rom[17098] = 16'hffff;
  rom[17099] = 16'hffff;
  rom[17100] = 16'hffff;
  rom[17101] = 16'hffff;
  rom[17102] = 16'hffff;
  rom[17103] = 16'hd67a;
  rom[17104] = 16'h2965;
  rom[17105] = 16'h10a2;
  rom[17106] = 16'h18a2;
  rom[17107] = 16'h2103;
  rom[17108] = 16'hbd96;
  rom[17109] = 16'hffff;
  rom[17110] = 16'hffff;
  rom[17111] = 16'hffff;
  rom[17112] = 16'hffff;
  rom[17113] = 16'hffff;
  rom[17114] = 16'hffff;
  rom[17115] = 16'hffdf;
  rom[17116] = 16'h9cd2;
  rom[17117] = 16'h2103;
  rom[17118] = 16'h18c2;
  rom[17119] = 16'h1082;
  rom[17120] = 16'h20c3;
  rom[17121] = 16'h18a2;
  rom[17122] = 16'h18c2;
  rom[17123] = 16'h18c2;
  rom[17124] = 16'h18c2;
  rom[17125] = 16'h10a2;
  rom[17126] = 16'h18e3;
  rom[17127] = 16'hce59;
  rom[17128] = 16'hffff;
  rom[17129] = 16'hffff;
  rom[17130] = 16'hffff;
  rom[17131] = 16'hffff;
  rom[17132] = 16'hffff;
  rom[17133] = 16'hffff;
  rom[17134] = 16'hffff;
  rom[17135] = 16'hffff;
  rom[17136] = 16'hffff;
  rom[17137] = 16'hffff;
  rom[17138] = 16'hffff;
  rom[17139] = 16'he6d9;
  rom[17140] = 16'h93aa;
  rom[17141] = 16'hcceb;
  rom[17142] = 16'hed8b;
  rom[17143] = 16'hf547;
  rom[17144] = 16'hfd68;
  rom[17145] = 16'hfd28;
  rom[17146] = 16'hfd4a;
  rom[17147] = 16'hf528;
  rom[17148] = 16'hfd49;
  rom[17149] = 16'hfd27;
  rom[17150] = 16'hfce7;
  rom[17151] = 16'hf529;
  rom[17152] = 16'hd50c;
  rom[17153] = 16'h7b28;
  rom[17154] = 16'hef1b;
  rom[17155] = 16'hffff;
  rom[17156] = 16'hffff;
  rom[17157] = 16'hffff;
  rom[17158] = 16'hffff;
  rom[17159] = 16'hffff;
  rom[17160] = 16'hffff;
  rom[17161] = 16'hffff;
  rom[17162] = 16'hffff;
  rom[17163] = 16'hffff;
  rom[17164] = 16'hffff;
  rom[17165] = 16'hffff;
  rom[17166] = 16'hffff;
  rom[17167] = 16'hffff;
  rom[17168] = 16'hffff;
  rom[17169] = 16'hffff;
  rom[17170] = 16'hffff;
  rom[17171] = 16'hffff;
  rom[17172] = 16'hffff;
  rom[17173] = 16'hffff;
  rom[17174] = 16'hffff;
  rom[17175] = 16'hffff;
  rom[17176] = 16'hffff;
  rom[17177] = 16'hffff;
  rom[17178] = 16'hffff;
  rom[17179] = 16'hffff;
  rom[17180] = 16'hffff;
  rom[17181] = 16'hffff;
  rom[17182] = 16'hffff;
  rom[17183] = 16'hffff;
  rom[17184] = 16'hffff;
  rom[17185] = 16'hffff;
  rom[17186] = 16'hffff;
  rom[17187] = 16'hffff;
  rom[17188] = 16'hffff;
  rom[17189] = 16'hffff;
  rom[17190] = 16'hffff;
  rom[17191] = 16'hffff;
  rom[17192] = 16'hffff;
  rom[17193] = 16'hffff;
  rom[17194] = 16'hffff;
  rom[17195] = 16'hffff;
  rom[17196] = 16'hffff;
  rom[17197] = 16'hffff;
  rom[17198] = 16'hffff;
  rom[17199] = 16'hffff;
  rom[17200] = 16'hffff;
  rom[17201] = 16'hffff;
  rom[17202] = 16'hffff;
  rom[17203] = 16'hffff;
  rom[17204] = 16'hffff;
  rom[17205] = 16'hffff;
  rom[17206] = 16'hffff;
  rom[17207] = 16'hffff;
  rom[17208] = 16'hffff;
  rom[17209] = 16'hffff;
  rom[17210] = 16'hffff;
  rom[17211] = 16'hffff;
  rom[17212] = 16'hffff;
  rom[17213] = 16'hffff;
  rom[17214] = 16'hffff;
  rom[17215] = 16'hffff;
  rom[17216] = 16'hffff;
  rom[17217] = 16'hffff;
  rom[17218] = 16'hffff;
  rom[17219] = 16'hffff;
  rom[17220] = 16'hffff;
  rom[17221] = 16'hffff;
  rom[17222] = 16'hffff;
  rom[17223] = 16'hffff;
  rom[17224] = 16'hffdf;
  rom[17225] = 16'hffff;
  rom[17226] = 16'hef9d;
  rom[17227] = 16'h7b89;
  rom[17228] = 16'hbd8b;
  rom[17229] = 16'hef0c;
  rom[17230] = 16'heee9;
  rom[17231] = 16'hff29;
  rom[17232] = 16'hf709;
  rom[17233] = 16'hff2a;
  rom[17234] = 16'hf729;
  rom[17235] = 16'hff28;
  rom[17236] = 16'hff08;
  rom[17237] = 16'hff28;
  rom[17238] = 16'hf708;
  rom[17239] = 16'hff28;
  rom[17240] = 16'hff08;
  rom[17241] = 16'hff28;
  rom[17242] = 16'hf708;
  rom[17243] = 16'hff28;
  rom[17244] = 16'hff08;
  rom[17245] = 16'hf709;
  rom[17246] = 16'hf70b;
  rom[17247] = 16'h9c23;
  rom[17248] = 16'h7a81;
  rom[17249] = 16'hdd09;
  rom[17250] = 16'hed48;
  rom[17251] = 16'hf54a;
  rom[17252] = 16'he529;
  rom[17253] = 16'hd52c;
  rom[17254] = 16'h7b48;
  rom[17255] = 16'hffdd;
  rom[17256] = 16'hfffe;
  rom[17257] = 16'hffff;
  rom[17258] = 16'hffff;
  rom[17259] = 16'hffff;
  rom[17260] = 16'hffff;
  rom[17261] = 16'hffff;
  rom[17262] = 16'hffff;
  rom[17263] = 16'hffff;
  rom[17264] = 16'hffdf;
  rom[17265] = 16'hffff;
  rom[17266] = 16'hffff;
  rom[17267] = 16'h842f;
  rom[17268] = 16'h20e3;
  rom[17269] = 16'h1082;
  rom[17270] = 16'h18a2;
  rom[17271] = 16'h18a2;
  rom[17272] = 16'h1081;
  rom[17273] = 16'h18a2;
  rom[17274] = 16'h18c3;
  rom[17275] = 16'h1082;
  rom[17276] = 16'h1082;
  rom[17277] = 16'h41e7;
  rom[17278] = 16'he6fb;
  rom[17279] = 16'hffbe;
  rom[17280] = 16'hffff;
  rom[17281] = 16'hffff;
  rom[17282] = 16'hffdf;
  rom[17283] = 16'hffff;
  rom[17284] = 16'hffff;
  rom[17285] = 16'hffdf;
  rom[17286] = 16'h7bcf;
  rom[17287] = 16'h18c2;
  rom[17288] = 16'h10a2;
  rom[17289] = 16'h2103;
  rom[17290] = 16'h8c50;
  rom[17291] = 16'hffff;
  rom[17292] = 16'hffff;
  rom[17293] = 16'hffff;
  rom[17294] = 16'hffff;
  rom[17295] = 16'hffff;
  rom[17296] = 16'hffff;
  rom[17297] = 16'hffff;
  rom[17298] = 16'hffff;
  rom[17299] = 16'hffff;
  rom[17300] = 16'hffff;
  rom[17301] = 16'hffff;
  rom[17302] = 16'hffff;
  rom[17303] = 16'hd6ba;
  rom[17304] = 16'h2945;
  rom[17305] = 16'h18e3;
  rom[17306] = 16'h10c2;
  rom[17307] = 16'h2945;
  rom[17308] = 16'had75;
  rom[17309] = 16'hffff;
  rom[17310] = 16'hffff;
  rom[17311] = 16'hffff;
  rom[17312] = 16'hffff;
  rom[17313] = 16'hffff;
  rom[17314] = 16'hffbe;
  rom[17315] = 16'hffff;
  rom[17316] = 16'h8c30;
  rom[17317] = 16'h18c3;
  rom[17318] = 16'h10a2;
  rom[17319] = 16'h18a2;
  rom[17320] = 16'h18a2;
  rom[17321] = 16'h18c2;
  rom[17322] = 16'h1081;
  rom[17323] = 16'h18a2;
  rom[17324] = 16'h18c2;
  rom[17325] = 16'h18c2;
  rom[17326] = 16'h20e3;
  rom[17327] = 16'hd69a;
  rom[17328] = 16'hffff;
  rom[17329] = 16'hffff;
  rom[17330] = 16'hffff;
  rom[17331] = 16'hffff;
  rom[17332] = 16'hffff;
  rom[17333] = 16'hffff;
  rom[17334] = 16'hffff;
  rom[17335] = 16'hffff;
  rom[17336] = 16'hffff;
  rom[17337] = 16'hffdf;
  rom[17338] = 16'hffde;
  rom[17339] = 16'hc592;
  rom[17340] = 16'h9387;
  rom[17341] = 16'he58d;
  rom[17342] = 16'hed69;
  rom[17343] = 16'hf588;
  rom[17344] = 16'hf547;
  rom[17345] = 16'hfd48;
  rom[17346] = 16'hf528;
  rom[17347] = 16'hf549;
  rom[17348] = 16'hfd28;
  rom[17349] = 16'hfd27;
  rom[17350] = 16'hf4e6;
  rom[17351] = 16'hf54a;
  rom[17352] = 16'hc4ec;
  rom[17353] = 16'h7b6a;
  rom[17354] = 16'hef5c;
  rom[17355] = 16'hffff;
  rom[17356] = 16'hffdf;
  rom[17357] = 16'hffff;
  rom[17358] = 16'hffff;
  rom[17359] = 16'hffff;
  rom[17360] = 16'hffff;
  rom[17361] = 16'hffff;
  rom[17362] = 16'hffff;
  rom[17363] = 16'hffff;
  rom[17364] = 16'hffff;
  rom[17365] = 16'hffff;
  rom[17366] = 16'hffff;
  rom[17367] = 16'hffff;
  rom[17368] = 16'hffff;
  rom[17369] = 16'hffff;
  rom[17370] = 16'hffff;
  rom[17371] = 16'hffff;
  rom[17372] = 16'hffff;
  rom[17373] = 16'hffff;
  rom[17374] = 16'hffff;
  rom[17375] = 16'hffff;
  rom[17376] = 16'hffff;
  rom[17377] = 16'hffff;
  rom[17378] = 16'hffff;
  rom[17379] = 16'hffff;
  rom[17380] = 16'hffff;
  rom[17381] = 16'hffff;
  rom[17382] = 16'hffff;
  rom[17383] = 16'hffff;
  rom[17384] = 16'hffff;
  rom[17385] = 16'hffff;
  rom[17386] = 16'hffff;
  rom[17387] = 16'hffff;
  rom[17388] = 16'hffff;
  rom[17389] = 16'hffff;
  rom[17390] = 16'hffff;
  rom[17391] = 16'hffff;
  rom[17392] = 16'hffff;
  rom[17393] = 16'hffff;
  rom[17394] = 16'hffff;
  rom[17395] = 16'hffff;
  rom[17396] = 16'hffff;
  rom[17397] = 16'hffff;
  rom[17398] = 16'hffff;
  rom[17399] = 16'hffff;
  rom[17400] = 16'hffff;
  rom[17401] = 16'hffff;
  rom[17402] = 16'hffff;
  rom[17403] = 16'hffff;
  rom[17404] = 16'hffff;
  rom[17405] = 16'hffff;
  rom[17406] = 16'hffff;
  rom[17407] = 16'hffff;
  rom[17408] = 16'hffff;
  rom[17409] = 16'hffff;
  rom[17410] = 16'hffff;
  rom[17411] = 16'hffff;
  rom[17412] = 16'hffff;
  rom[17413] = 16'hffff;
  rom[17414] = 16'hffff;
  rom[17415] = 16'hffff;
  rom[17416] = 16'hffff;
  rom[17417] = 16'hffff;
  rom[17418] = 16'hffff;
  rom[17419] = 16'hffff;
  rom[17420] = 16'hffff;
  rom[17421] = 16'hffff;
  rom[17422] = 16'hffff;
  rom[17423] = 16'hffff;
  rom[17424] = 16'hffff;
  rom[17425] = 16'hffff;
  rom[17426] = 16'hef7c;
  rom[17427] = 16'h62e5;
  rom[17428] = 16'hd64d;
  rom[17429] = 16'hf70b;
  rom[17430] = 16'hff2a;
  rom[17431] = 16'hff49;
  rom[17432] = 16'hff29;
  rom[17433] = 16'hf729;
  rom[17434] = 16'hff29;
  rom[17435] = 16'hff28;
  rom[17436] = 16'hff29;
  rom[17437] = 16'hff29;
  rom[17438] = 16'hff29;
  rom[17439] = 16'hff28;
  rom[17440] = 16'hff29;
  rom[17441] = 16'hff28;
  rom[17442] = 16'hff29;
  rom[17443] = 16'hff28;
  rom[17444] = 16'hff29;
  rom[17445] = 16'hf74a;
  rom[17446] = 16'hf70b;
  rom[17447] = 16'hddea;
  rom[17448] = 16'h6a01;
  rom[17449] = 16'hd4a9;
  rom[17450] = 16'hed28;
  rom[17451] = 16'hf549;
  rom[17452] = 16'hf56a;
  rom[17453] = 16'hd50a;
  rom[17454] = 16'h9347;
  rom[17455] = 16'hc573;
  rom[17456] = 16'hfffe;
  rom[17457] = 16'hffff;
  rom[17458] = 16'hffff;
  rom[17459] = 16'hffff;
  rom[17460] = 16'hffff;
  rom[17461] = 16'hffff;
  rom[17462] = 16'hffff;
  rom[17463] = 16'hffff;
  rom[17464] = 16'hffff;
  rom[17465] = 16'hffff;
  rom[17466] = 16'hffff;
  rom[17467] = 16'hbdd7;
  rom[17468] = 16'h20e3;
  rom[17469] = 16'h1082;
  rom[17470] = 16'h2103;
  rom[17471] = 16'h10a2;
  rom[17472] = 16'h20e3;
  rom[17473] = 16'h18a2;
  rom[17474] = 16'h20c3;
  rom[17475] = 16'h18a2;
  rom[17476] = 16'h18c3;
  rom[17477] = 16'h2924;
  rom[17478] = 16'hce58;
  rom[17479] = 16'hffdf;
  rom[17480] = 16'hffff;
  rom[17481] = 16'hffdf;
  rom[17482] = 16'hffff;
  rom[17483] = 16'hffdf;
  rom[17484] = 16'hffff;
  rom[17485] = 16'hd69a;
  rom[17486] = 16'h4207;
  rom[17487] = 16'h1081;
  rom[17488] = 16'h2104;
  rom[17489] = 16'h18c2;
  rom[17490] = 16'hc5f7;
  rom[17491] = 16'hffff;
  rom[17492] = 16'hffff;
  rom[17493] = 16'hffff;
  rom[17494] = 16'hffff;
  rom[17495] = 16'hffff;
  rom[17496] = 16'hffff;
  rom[17497] = 16'hffff;
  rom[17498] = 16'hffff;
  rom[17499] = 16'hffff;
  rom[17500] = 16'hffff;
  rom[17501] = 16'hffff;
  rom[17502] = 16'hffff;
  rom[17503] = 16'hef5c;
  rom[17504] = 16'h5269;
  rom[17505] = 16'h18c2;
  rom[17506] = 16'h18e3;
  rom[17507] = 16'h18e2;
  rom[17508] = 16'h8c51;
  rom[17509] = 16'hf79e;
  rom[17510] = 16'hffff;
  rom[17511] = 16'hffff;
  rom[17512] = 16'hffff;
  rom[17513] = 16'hffff;
  rom[17514] = 16'hffdf;
  rom[17515] = 16'hef3c;
  rom[17516] = 16'h62eb;
  rom[17517] = 16'h18c2;
  rom[17518] = 16'h18c2;
  rom[17519] = 16'h18c2;
  rom[17520] = 16'h18a3;
  rom[17521] = 16'h18a2;
  rom[17522] = 16'h20e3;
  rom[17523] = 16'h10c2;
  rom[17524] = 16'h18e3;
  rom[17525] = 16'h10c2;
  rom[17526] = 16'h4a29;
  rom[17527] = 16'he6fb;
  rom[17528] = 16'hffff;
  rom[17529] = 16'hffff;
  rom[17530] = 16'hffff;
  rom[17531] = 16'hffff;
  rom[17532] = 16'hffff;
  rom[17533] = 16'hffff;
  rom[17534] = 16'hffff;
  rom[17535] = 16'hffff;
  rom[17536] = 16'hffff;
  rom[17537] = 16'hffff;
  rom[17538] = 16'hffdc;
  rom[17539] = 16'h93ea;
  rom[17540] = 16'hc48a;
  rom[17541] = 16'he54a;
  rom[17542] = 16'hf58a;
  rom[17543] = 16'hf568;
  rom[17544] = 16'hfd68;
  rom[17545] = 16'hfd28;
  rom[17546] = 16'hfd28;
  rom[17547] = 16'hfd29;
  rom[17548] = 16'hfd49;
  rom[17549] = 16'hfd07;
  rom[17550] = 16'hfd07;
  rom[17551] = 16'hed4a;
  rom[17552] = 16'ha40a;
  rom[17553] = 16'h9c6e;
  rom[17554] = 16'hf79d;
  rom[17555] = 16'hffdf;
  rom[17556] = 16'hffff;
  rom[17557] = 16'hffff;
  rom[17558] = 16'hffff;
  rom[17559] = 16'hffff;
  rom[17560] = 16'hffff;
  rom[17561] = 16'hffff;
  rom[17562] = 16'hffff;
  rom[17563] = 16'hffff;
  rom[17564] = 16'hffff;
  rom[17565] = 16'hffff;
  rom[17566] = 16'hffff;
  rom[17567] = 16'hffff;
  rom[17568] = 16'hffff;
  rom[17569] = 16'hffff;
  rom[17570] = 16'hffff;
  rom[17571] = 16'hffff;
  rom[17572] = 16'hffff;
  rom[17573] = 16'hffff;
  rom[17574] = 16'hffff;
  rom[17575] = 16'hffff;
  rom[17576] = 16'hffff;
  rom[17577] = 16'hffff;
  rom[17578] = 16'hffff;
  rom[17579] = 16'hffff;
  rom[17580] = 16'hffff;
  rom[17581] = 16'hffff;
  rom[17582] = 16'hffff;
  rom[17583] = 16'hffff;
  rom[17584] = 16'hffff;
  rom[17585] = 16'hffff;
  rom[17586] = 16'hffff;
  rom[17587] = 16'hffff;
  rom[17588] = 16'hffff;
  rom[17589] = 16'hffff;
  rom[17590] = 16'hffff;
  rom[17591] = 16'hffff;
  rom[17592] = 16'hffff;
  rom[17593] = 16'hffff;
  rom[17594] = 16'hffff;
  rom[17595] = 16'hffff;
  rom[17596] = 16'hffff;
  rom[17597] = 16'hffff;
  rom[17598] = 16'hffff;
  rom[17599] = 16'hffff;
  rom[17600] = 16'hffff;
  rom[17601] = 16'hffff;
  rom[17602] = 16'hffff;
  rom[17603] = 16'hffff;
  rom[17604] = 16'hffff;
  rom[17605] = 16'hffff;
  rom[17606] = 16'hffff;
  rom[17607] = 16'hffff;
  rom[17608] = 16'hffff;
  rom[17609] = 16'hffff;
  rom[17610] = 16'hffff;
  rom[17611] = 16'hffff;
  rom[17612] = 16'hffff;
  rom[17613] = 16'hffff;
  rom[17614] = 16'hffff;
  rom[17615] = 16'hffff;
  rom[17616] = 16'hffff;
  rom[17617] = 16'hffff;
  rom[17618] = 16'hffff;
  rom[17619] = 16'hffff;
  rom[17620] = 16'hffff;
  rom[17621] = 16'hffff;
  rom[17622] = 16'hffff;
  rom[17623] = 16'hffff;
  rom[17624] = 16'hffdf;
  rom[17625] = 16'hffff;
  rom[17626] = 16'hef5a;
  rom[17627] = 16'h62e3;
  rom[17628] = 16'hd60a;
  rom[17629] = 16'hf70a;
  rom[17630] = 16'hf6e8;
  rom[17631] = 16'hff29;
  rom[17632] = 16'hf728;
  rom[17633] = 16'hff28;
  rom[17634] = 16'hff08;
  rom[17635] = 16'hff29;
  rom[17636] = 16'hf709;
  rom[17637] = 16'hff29;
  rom[17638] = 16'hff09;
  rom[17639] = 16'hff29;
  rom[17640] = 16'hf708;
  rom[17641] = 16'hff28;
  rom[17642] = 16'hff08;
  rom[17643] = 16'hff28;
  rom[17644] = 16'hf708;
  rom[17645] = 16'hf709;
  rom[17646] = 16'hf72b;
  rom[17647] = 16'hf6ed;
  rom[17648] = 16'h7240;
  rom[17649] = 16'hb406;
  rom[17650] = 16'hf5aa;
  rom[17651] = 16'hf549;
  rom[17652] = 16'hed28;
  rom[17653] = 16'hf58b;
  rom[17654] = 16'hbc49;
  rom[17655] = 16'h8328;
  rom[17656] = 16'hf79c;
  rom[17657] = 16'hffff;
  rom[17658] = 16'hffff;
  rom[17659] = 16'hffff;
  rom[17660] = 16'hffff;
  rom[17661] = 16'hffff;
  rom[17662] = 16'hffff;
  rom[17663] = 16'hffff;
  rom[17664] = 16'hffbe;
  rom[17665] = 16'hffff;
  rom[17666] = 16'hffff;
  rom[17667] = 16'hde9a;
  rom[17668] = 16'h39a6;
  rom[17669] = 16'h18a2;
  rom[17670] = 16'h18a2;
  rom[17671] = 16'h18a2;
  rom[17672] = 16'h1082;
  rom[17673] = 16'h18c2;
  rom[17674] = 16'h1061;
  rom[17675] = 16'h20c3;
  rom[17676] = 16'h2103;
  rom[17677] = 16'h1061;
  rom[17678] = 16'h5aaa;
  rom[17679] = 16'hd659;
  rom[17680] = 16'hffdf;
  rom[17681] = 16'hffff;
  rom[17682] = 16'hffdf;
  rom[17683] = 16'hffff;
  rom[17684] = 16'hf77d;
  rom[17685] = 16'h83ef;
  rom[17686] = 16'h10a2;
  rom[17687] = 16'h18c3;
  rom[17688] = 16'h2104;
  rom[17689] = 16'h31a6;
  rom[17690] = 16'he71c;
  rom[17691] = 16'hffdf;
  rom[17692] = 16'hffff;
  rom[17693] = 16'hffff;
  rom[17694] = 16'hffff;
  rom[17695] = 16'hffff;
  rom[17696] = 16'hffff;
  rom[17697] = 16'hffff;
  rom[17698] = 16'hffff;
  rom[17699] = 16'hffff;
  rom[17700] = 16'hffff;
  rom[17701] = 16'hffff;
  rom[17702] = 16'hffff;
  rom[17703] = 16'hffbf;
  rom[17704] = 16'h7bce;
  rom[17705] = 16'h18c3;
  rom[17706] = 16'h10a1;
  rom[17707] = 16'h10a2;
  rom[17708] = 16'h39c6;
  rom[17709] = 16'hbdd6;
  rom[17710] = 16'hffff;
  rom[17711] = 16'hffff;
  rom[17712] = 16'hffde;
  rom[17713] = 16'hffff;
  rom[17714] = 16'hffdf;
  rom[17715] = 16'ha514;
  rom[17716] = 16'h2123;
  rom[17717] = 16'h18a2;
  rom[17718] = 16'h18a2;
  rom[17719] = 16'h18a2;
  rom[17720] = 16'h1082;
  rom[17721] = 16'h18c2;
  rom[17722] = 16'h18a2;
  rom[17723] = 16'h18c2;
  rom[17724] = 16'h10c2;
  rom[17725] = 16'h18c2;
  rom[17726] = 16'h9451;
  rom[17727] = 16'hffbf;
  rom[17728] = 16'hffff;
  rom[17729] = 16'hffff;
  rom[17730] = 16'hffff;
  rom[17731] = 16'hffff;
  rom[17732] = 16'hffff;
  rom[17733] = 16'hffff;
  rom[17734] = 16'hffff;
  rom[17735] = 16'hffff;
  rom[17736] = 16'hffdf;
  rom[17737] = 16'hfffe;
  rom[17738] = 16'hd634;
  rom[17739] = 16'h8b26;
  rom[17740] = 16'hdd2b;
  rom[17741] = 16'hed4a;
  rom[17742] = 16'hf569;
  rom[17743] = 16'hf568;
  rom[17744] = 16'hf547;
  rom[17745] = 16'hfd47;
  rom[17746] = 16'hfd27;
  rom[17747] = 16'hf529;
  rom[17748] = 16'hfd08;
  rom[17749] = 16'hfd48;
  rom[17750] = 16'hf4e7;
  rom[17751] = 16'he54b;
  rom[17752] = 16'h8347;
  rom[17753] = 16'ha532;
  rom[17754] = 16'hef7d;
  rom[17755] = 16'hffff;
  rom[17756] = 16'hffff;
  rom[17757] = 16'hffff;
  rom[17758] = 16'hffff;
  rom[17759] = 16'hffff;
  rom[17760] = 16'hffff;
  rom[17761] = 16'hffff;
  rom[17762] = 16'hffff;
  rom[17763] = 16'hffff;
  rom[17764] = 16'hffff;
  rom[17765] = 16'hffff;
  rom[17766] = 16'hffff;
  rom[17767] = 16'hffff;
  rom[17768] = 16'hffff;
  rom[17769] = 16'hffff;
  rom[17770] = 16'hffff;
  rom[17771] = 16'hffff;
  rom[17772] = 16'hffff;
  rom[17773] = 16'hffff;
  rom[17774] = 16'hffff;
  rom[17775] = 16'hffff;
  rom[17776] = 16'hffff;
  rom[17777] = 16'hffff;
  rom[17778] = 16'hffff;
  rom[17779] = 16'hffff;
  rom[17780] = 16'hffff;
  rom[17781] = 16'hffff;
  rom[17782] = 16'hffff;
  rom[17783] = 16'hffff;
  rom[17784] = 16'hffff;
  rom[17785] = 16'hffff;
  rom[17786] = 16'hffff;
  rom[17787] = 16'hffff;
  rom[17788] = 16'hffff;
  rom[17789] = 16'hffff;
  rom[17790] = 16'hffff;
  rom[17791] = 16'hffff;
  rom[17792] = 16'hffff;
  rom[17793] = 16'hffff;
  rom[17794] = 16'hffff;
  rom[17795] = 16'hffff;
  rom[17796] = 16'hffff;
  rom[17797] = 16'hffff;
  rom[17798] = 16'hffff;
  rom[17799] = 16'hffff;
  rom[17800] = 16'hffff;
  rom[17801] = 16'hffff;
  rom[17802] = 16'hffff;
  rom[17803] = 16'hffff;
  rom[17804] = 16'hffff;
  rom[17805] = 16'hffff;
  rom[17806] = 16'hffff;
  rom[17807] = 16'hffff;
  rom[17808] = 16'hffff;
  rom[17809] = 16'hffff;
  rom[17810] = 16'hffff;
  rom[17811] = 16'hffff;
  rom[17812] = 16'hffff;
  rom[17813] = 16'hffff;
  rom[17814] = 16'hffff;
  rom[17815] = 16'hffff;
  rom[17816] = 16'hffff;
  rom[17817] = 16'hffff;
  rom[17818] = 16'hffff;
  rom[17819] = 16'hffff;
  rom[17820] = 16'hffff;
  rom[17821] = 16'hffff;
  rom[17822] = 16'hffff;
  rom[17823] = 16'hffff;
  rom[17824] = 16'hffff;
  rom[17825] = 16'hffff;
  rom[17826] = 16'hf77b;
  rom[17827] = 16'h5aa1;
  rom[17828] = 16'hde6b;
  rom[17829] = 16'hf70a;
  rom[17830] = 16'hff2a;
  rom[17831] = 16'hff29;
  rom[17832] = 16'hff29;
  rom[17833] = 16'hf727;
  rom[17834] = 16'hff29;
  rom[17835] = 16'hff29;
  rom[17836] = 16'hff2a;
  rom[17837] = 16'hff29;
  rom[17838] = 16'hff2a;
  rom[17839] = 16'hff29;
  rom[17840] = 16'hff2a;
  rom[17841] = 16'hff28;
  rom[17842] = 16'hff29;
  rom[17843] = 16'hff28;
  rom[17844] = 16'hff29;
  rom[17845] = 16'hf749;
  rom[17846] = 16'hff2b;
  rom[17847] = 16'hcd88;
  rom[17848] = 16'h6a22;
  rom[17849] = 16'hcc89;
  rom[17850] = 16'hf58b;
  rom[17851] = 16'hfd69;
  rom[17852] = 16'hf507;
  rom[17853] = 16'hfd8a;
  rom[17854] = 16'hdceb;
  rom[17855] = 16'h9348;
  rom[17856] = 16'hc574;
  rom[17857] = 16'hffff;
  rom[17858] = 16'hffff;
  rom[17859] = 16'hffff;
  rom[17860] = 16'hffff;
  rom[17861] = 16'hffff;
  rom[17862] = 16'hffff;
  rom[17863] = 16'hffff;
  rom[17864] = 16'hffff;
  rom[17865] = 16'hffff;
  rom[17866] = 16'hffff;
  rom[17867] = 16'hf79e;
  rom[17868] = 16'h7bae;
  rom[17869] = 16'h18a3;
  rom[17870] = 16'h18a3;
  rom[17871] = 16'h18c3;
  rom[17872] = 16'h18a2;
  rom[17873] = 16'h18a2;
  rom[17874] = 16'h2904;
  rom[17875] = 16'h18a2;
  rom[17876] = 16'h20c2;
  rom[17877] = 16'h18c2;
  rom[17878] = 16'h1882;
  rom[17879] = 16'h52aa;
  rom[17880] = 16'had34;
  rom[17881] = 16'hce59;
  rom[17882] = 16'hdeba;
  rom[17883] = 16'hb575;
  rom[17884] = 16'h6b2c;
  rom[17885] = 16'h2123;
  rom[17886] = 16'h18c3;
  rom[17887] = 16'h18e3;
  rom[17888] = 16'h1061;
  rom[17889] = 16'h73ae;
  rom[17890] = 16'hff9e;
  rom[17891] = 16'hffff;
  rom[17892] = 16'hffff;
  rom[17893] = 16'hffff;
  rom[17894] = 16'hffff;
  rom[17895] = 16'hffff;
  rom[17896] = 16'hffff;
  rom[17897] = 16'hffff;
  rom[17898] = 16'hffff;
  rom[17899] = 16'hffff;
  rom[17900] = 16'hffff;
  rom[17901] = 16'hffff;
  rom[17902] = 16'hffff;
  rom[17903] = 16'hffff;
  rom[17904] = 16'hd679;
  rom[17905] = 16'h18c3;
  rom[17906] = 16'h20c3;
  rom[17907] = 16'h20e3;
  rom[17908] = 16'h18a2;
  rom[17909] = 16'h4228;
  rom[17910] = 16'h9451;
  rom[17911] = 16'hce18;
  rom[17912] = 16'hdebb;
  rom[17913] = 16'hc618;
  rom[17914] = 16'h83ef;
  rom[17915] = 16'h39a6;
  rom[17916] = 16'h18e3;
  rom[17917] = 16'h18a2;
  rom[17918] = 16'h18c2;
  rom[17919] = 16'h18a2;
  rom[17920] = 16'h20e3;
  rom[17921] = 16'h18c2;
  rom[17922] = 16'h18a2;
  rom[17923] = 16'h18c2;
  rom[17924] = 16'h18c2;
  rom[17925] = 16'h39e7;
  rom[17926] = 16'hd69a;
  rom[17927] = 16'hffff;
  rom[17928] = 16'hffff;
  rom[17929] = 16'hffff;
  rom[17930] = 16'hffff;
  rom[17931] = 16'hffff;
  rom[17932] = 16'hffff;
  rom[17933] = 16'hffff;
  rom[17934] = 16'hffff;
  rom[17935] = 16'hffff;
  rom[17936] = 16'hffff;
  rom[17937] = 16'hef3a;
  rom[17938] = 16'h8388;
  rom[17939] = 16'hac28;
  rom[17940] = 16'hed4b;
  rom[17941] = 16'hf56a;
  rom[17942] = 16'hfd49;
  rom[17943] = 16'hf548;
  rom[17944] = 16'hfd47;
  rom[17945] = 16'hfd27;
  rom[17946] = 16'hfd28;
  rom[17947] = 16'hfd49;
  rom[17948] = 16'hfd09;
  rom[17949] = 16'hfd08;
  rom[17950] = 16'hfd69;
  rom[17951] = 16'hdcea;
  rom[17952] = 16'h7b48;
  rom[17953] = 16'hbdf6;
  rom[17954] = 16'hffff;
  rom[17955] = 16'hffff;
  rom[17956] = 16'hffdf;
  rom[17957] = 16'hffff;
  rom[17958] = 16'hffff;
  rom[17959] = 16'hffff;
  rom[17960] = 16'hffff;
  rom[17961] = 16'hffff;
  rom[17962] = 16'hffff;
  rom[17963] = 16'hffff;
  rom[17964] = 16'hffff;
  rom[17965] = 16'hffff;
  rom[17966] = 16'hffff;
  rom[17967] = 16'hffff;
  rom[17968] = 16'hffff;
  rom[17969] = 16'hffff;
  rom[17970] = 16'hffff;
  rom[17971] = 16'hffff;
  rom[17972] = 16'hffff;
  rom[17973] = 16'hffff;
  rom[17974] = 16'hffff;
  rom[17975] = 16'hffff;
  rom[17976] = 16'hffff;
  rom[17977] = 16'hffff;
  rom[17978] = 16'hffff;
  rom[17979] = 16'hffff;
  rom[17980] = 16'hffff;
  rom[17981] = 16'hffff;
  rom[17982] = 16'hffff;
  rom[17983] = 16'hffff;
  rom[17984] = 16'hffff;
  rom[17985] = 16'hffff;
  rom[17986] = 16'hffff;
  rom[17987] = 16'hffff;
  rom[17988] = 16'hffff;
  rom[17989] = 16'hffff;
  rom[17990] = 16'hffff;
  rom[17991] = 16'hffff;
  rom[17992] = 16'hffff;
  rom[17993] = 16'hffff;
  rom[17994] = 16'hffff;
  rom[17995] = 16'hffff;
  rom[17996] = 16'hffff;
  rom[17997] = 16'hffff;
  rom[17998] = 16'hffff;
  rom[17999] = 16'hffff;
  rom[18000] = 16'hffff;
  rom[18001] = 16'hffff;
  rom[18002] = 16'hffff;
  rom[18003] = 16'hffff;
  rom[18004] = 16'hffff;
  rom[18005] = 16'hffff;
  rom[18006] = 16'hffff;
  rom[18007] = 16'hffff;
  rom[18008] = 16'hffff;
  rom[18009] = 16'hffff;
  rom[18010] = 16'hffff;
  rom[18011] = 16'hffff;
  rom[18012] = 16'hffff;
  rom[18013] = 16'hffff;
  rom[18014] = 16'hffff;
  rom[18015] = 16'hffff;
  rom[18016] = 16'hffff;
  rom[18017] = 16'hffff;
  rom[18018] = 16'hffff;
  rom[18019] = 16'hffff;
  rom[18020] = 16'hffff;
  rom[18021] = 16'hffff;
  rom[18022] = 16'hffff;
  rom[18023] = 16'hffff;
  rom[18024] = 16'hffdf;
  rom[18025] = 16'hffff;
  rom[18026] = 16'he739;
  rom[18027] = 16'h5a81;
  rom[18028] = 16'hde6a;
  rom[18029] = 16'hff0a;
  rom[18030] = 16'hf6e9;
  rom[18031] = 16'hff0a;
  rom[18032] = 16'hff09;
  rom[18033] = 16'hff28;
  rom[18034] = 16'hf708;
  rom[18035] = 16'hff29;
  rom[18036] = 16'hff09;
  rom[18037] = 16'hff29;
  rom[18038] = 16'hf709;
  rom[18039] = 16'hff29;
  rom[18040] = 16'hff08;
  rom[18041] = 16'hff28;
  rom[18042] = 16'hf708;
  rom[18043] = 16'hff28;
  rom[18044] = 16'hf708;
  rom[18045] = 16'hf749;
  rom[18046] = 16'hf72a;
  rom[18047] = 16'hbce4;
  rom[18048] = 16'h61e1;
  rom[18049] = 16'hccea;
  rom[18050] = 16'he549;
  rom[18051] = 16'hf548;
  rom[18052] = 16'hfd27;
  rom[18053] = 16'hfce8;
  rom[18054] = 16'hf52b;
  rom[18055] = 16'hbc6b;
  rom[18056] = 16'h8baa;
  rom[18057] = 16'hf75b;
  rom[18058] = 16'hffff;
  rom[18059] = 16'hffff;
  rom[18060] = 16'hffff;
  rom[18061] = 16'hffff;
  rom[18062] = 16'hffff;
  rom[18063] = 16'hffff;
  rom[18064] = 16'hffdf;
  rom[18065] = 16'hffff;
  rom[18066] = 16'hffff;
  rom[18067] = 16'hffff;
  rom[18068] = 16'hc618;
  rom[18069] = 16'h2965;
  rom[18070] = 16'h1081;
  rom[18071] = 16'h18e3;
  rom[18072] = 16'h18a2;
  rom[18073] = 16'h18c3;
  rom[18074] = 16'h1081;
  rom[18075] = 16'h20e3;
  rom[18076] = 16'h1082;
  rom[18077] = 16'h18a2;
  rom[18078] = 16'h1081;
  rom[18079] = 16'h18e3;
  rom[18080] = 16'h18c2;
  rom[18081] = 16'h3986;
  rom[18082] = 16'h3185;
  rom[18083] = 16'h2144;
  rom[18084] = 16'h10a2;
  rom[18085] = 16'h18c3;
  rom[18086] = 16'h10a2;
  rom[18087] = 16'h10a2;
  rom[18088] = 16'h3145;
  rom[18089] = 16'hce39;
  rom[18090] = 16'hffff;
  rom[18091] = 16'hffff;
  rom[18092] = 16'hffff;
  rom[18093] = 16'hffff;
  rom[18094] = 16'hffff;
  rom[18095] = 16'hffff;
  rom[18096] = 16'hffff;
  rom[18097] = 16'hffff;
  rom[18098] = 16'hffff;
  rom[18099] = 16'hffff;
  rom[18100] = 16'hffff;
  rom[18101] = 16'hffff;
  rom[18102] = 16'hffff;
  rom[18103] = 16'hffff;
  rom[18104] = 16'hffdf;
  rom[18105] = 16'h83ef;
  rom[18106] = 16'h10a2;
  rom[18107] = 16'h18e3;
  rom[18108] = 16'h18c2;
  rom[18109] = 16'h18c3;
  rom[18110] = 16'h18c2;
  rom[18111] = 16'h31a6;
  rom[18112] = 16'h3186;
  rom[18113] = 16'h3165;
  rom[18114] = 16'h18c2;
  rom[18115] = 16'h18a2;
  rom[18116] = 16'h10a1;
  rom[18117] = 16'h18c2;
  rom[18118] = 16'h10a1;
  rom[18119] = 16'h18a2;
  rom[18120] = 16'h18a1;
  rom[18121] = 16'h18a2;
  rom[18122] = 16'h18a2;
  rom[18123] = 16'h1081;
  rom[18124] = 16'h18c1;
  rom[18125] = 16'h7bcf;
  rom[18126] = 16'hf7be;
  rom[18127] = 16'hffff;
  rom[18128] = 16'hffdf;
  rom[18129] = 16'hffff;
  rom[18130] = 16'hffff;
  rom[18131] = 16'hffff;
  rom[18132] = 16'hffff;
  rom[18133] = 16'hffff;
  rom[18134] = 16'hffff;
  rom[18135] = 16'hffff;
  rom[18136] = 16'hffff;
  rom[18137] = 16'hb530;
  rom[18138] = 16'h7b45;
  rom[18139] = 16'hd50a;
  rom[18140] = 16'hfd6b;
  rom[18141] = 16'hfd08;
  rom[18142] = 16'hfd28;
  rom[18143] = 16'hf527;
  rom[18144] = 16'hf547;
  rom[18145] = 16'hfd47;
  rom[18146] = 16'hf527;
  rom[18147] = 16'hf529;
  rom[18148] = 16'hfd08;
  rom[18149] = 16'hfce8;
  rom[18150] = 16'hfd6b;
  rom[18151] = 16'hc449;
  rom[18152] = 16'h8369;
  rom[18153] = 16'he71c;
  rom[18154] = 16'hffff;
  rom[18155] = 16'hffff;
  rom[18156] = 16'hffff;
  rom[18157] = 16'hffff;
  rom[18158] = 16'hffff;
  rom[18159] = 16'hffff;
  rom[18160] = 16'hffff;
  rom[18161] = 16'hffff;
  rom[18162] = 16'hffff;
  rom[18163] = 16'hffff;
  rom[18164] = 16'hffff;
  rom[18165] = 16'hffff;
  rom[18166] = 16'hffff;
  rom[18167] = 16'hffff;
  rom[18168] = 16'hffff;
  rom[18169] = 16'hffff;
  rom[18170] = 16'hffff;
  rom[18171] = 16'hffff;
  rom[18172] = 16'hffff;
  rom[18173] = 16'hffff;
  rom[18174] = 16'hffff;
  rom[18175] = 16'hffff;
  rom[18176] = 16'hffff;
  rom[18177] = 16'hffff;
  rom[18178] = 16'hffff;
  rom[18179] = 16'hffff;
  rom[18180] = 16'hffff;
  rom[18181] = 16'hffff;
  rom[18182] = 16'hffff;
  rom[18183] = 16'hffff;
  rom[18184] = 16'hffff;
  rom[18185] = 16'hffff;
  rom[18186] = 16'hffff;
  rom[18187] = 16'hffff;
  rom[18188] = 16'hffff;
  rom[18189] = 16'hffff;
  rom[18190] = 16'hffff;
  rom[18191] = 16'hffff;
  rom[18192] = 16'hffff;
  rom[18193] = 16'hffff;
  rom[18194] = 16'hffff;
  rom[18195] = 16'hffff;
  rom[18196] = 16'hffff;
  rom[18197] = 16'hffff;
  rom[18198] = 16'hffff;
  rom[18199] = 16'hffff;
  rom[18200] = 16'hffff;
  rom[18201] = 16'hffff;
  rom[18202] = 16'hffff;
  rom[18203] = 16'hffff;
  rom[18204] = 16'hffff;
  rom[18205] = 16'hffff;
  rom[18206] = 16'hffff;
  rom[18207] = 16'hffff;
  rom[18208] = 16'hffff;
  rom[18209] = 16'hffff;
  rom[18210] = 16'hffff;
  rom[18211] = 16'hffff;
  rom[18212] = 16'hffff;
  rom[18213] = 16'hffff;
  rom[18214] = 16'hffff;
  rom[18215] = 16'hffff;
  rom[18216] = 16'hffff;
  rom[18217] = 16'hffff;
  rom[18218] = 16'hffff;
  rom[18219] = 16'hffff;
  rom[18220] = 16'hffff;
  rom[18221] = 16'hffff;
  rom[18222] = 16'hffff;
  rom[18223] = 16'hffff;
  rom[18224] = 16'hffff;
  rom[18225] = 16'hffff;
  rom[18226] = 16'hef3a;
  rom[18227] = 16'h5ac2;
  rom[18228] = 16'hd62a;
  rom[18229] = 16'hff2a;
  rom[18230] = 16'hff0a;
  rom[18231] = 16'hff0a;
  rom[18232] = 16'hff2a;
  rom[18233] = 16'hf709;
  rom[18234] = 16'hff2a;
  rom[18235] = 16'hff29;
  rom[18236] = 16'hff29;
  rom[18237] = 16'hff29;
  rom[18238] = 16'hff29;
  rom[18239] = 16'hff29;
  rom[18240] = 16'hff29;
  rom[18241] = 16'hff28;
  rom[18242] = 16'hff29;
  rom[18243] = 16'hff28;
  rom[18244] = 16'hff29;
  rom[18245] = 16'hf749;
  rom[18246] = 16'hf72a;
  rom[18247] = 16'hde27;
  rom[18248] = 16'h82c1;
  rom[18249] = 16'habe7;
  rom[18250] = 16'he56b;
  rom[18251] = 16'hf568;
  rom[18252] = 16'hfd48;
  rom[18253] = 16'hfcc7;
  rom[18254] = 16'hfd6b;
  rom[18255] = 16'hd4ea;
  rom[18256] = 16'h9be9;
  rom[18257] = 16'h9c8f;
  rom[18258] = 16'hff7d;
  rom[18259] = 16'hffdf;
  rom[18260] = 16'hffff;
  rom[18261] = 16'hffff;
  rom[18262] = 16'hffff;
  rom[18263] = 16'hfffe;
  rom[18264] = 16'hffff;
  rom[18265] = 16'hffff;
  rom[18266] = 16'hffff;
  rom[18267] = 16'hffff;
  rom[18268] = 16'hffbe;
  rom[18269] = 16'h9cb2;
  rom[18270] = 16'h3166;
  rom[18271] = 16'h10a2;
  rom[18272] = 16'h18a2;
  rom[18273] = 16'h20c3;
  rom[18274] = 16'h1882;
  rom[18275] = 16'h18a2;
  rom[18276] = 16'h3145;
  rom[18277] = 16'h1082;
  rom[18278] = 16'h20e4;
  rom[18279] = 16'h18c3;
  rom[18280] = 16'h18a2;
  rom[18281] = 16'h2944;
  rom[18282] = 16'h18c2;
  rom[18283] = 16'h10c2;
  rom[18284] = 16'h18c2;
  rom[18285] = 16'h18a2;
  rom[18286] = 16'h18c2;
  rom[18287] = 16'h2944;
  rom[18288] = 16'had34;
  rom[18289] = 16'hffff;
  rom[18290] = 16'hffff;
  rom[18291] = 16'hffff;
  rom[18292] = 16'hffff;
  rom[18293] = 16'hffff;
  rom[18294] = 16'hffff;
  rom[18295] = 16'hffff;
  rom[18296] = 16'hffff;
  rom[18297] = 16'hffff;
  rom[18298] = 16'hffff;
  rom[18299] = 16'hffff;
  rom[18300] = 16'hffff;
  rom[18301] = 16'hffff;
  rom[18302] = 16'hffff;
  rom[18303] = 16'hffff;
  rom[18304] = 16'hffff;
  rom[18305] = 16'hf77e;
  rom[18306] = 16'h5aaa;
  rom[18307] = 16'h18c3;
  rom[18308] = 16'h18c3;
  rom[18309] = 16'h18a2;
  rom[18310] = 16'h18c3;
  rom[18311] = 16'h18c2;
  rom[18312] = 16'h18c3;
  rom[18313] = 16'h20e3;
  rom[18314] = 16'h20c3;
  rom[18315] = 16'h18c2;
  rom[18316] = 16'h20c3;
  rom[18317] = 16'h18a2;
  rom[18318] = 16'h20e3;
  rom[18319] = 16'h18a2;
  rom[18320] = 16'h18a2;
  rom[18321] = 16'h18a2;
  rom[18322] = 16'h18a2;
  rom[18323] = 16'h20c2;
  rom[18324] = 16'h5a89;
  rom[18325] = 16'hd679;
  rom[18326] = 16'hffff;
  rom[18327] = 16'hffff;
  rom[18328] = 16'hffff;
  rom[18329] = 16'hffff;
  rom[18330] = 16'hffff;
  rom[18331] = 16'hffff;
  rom[18332] = 16'hffff;
  rom[18333] = 16'hffff;
  rom[18334] = 16'hffff;
  rom[18335] = 16'hff9e;
  rom[18336] = 16'he6b9;
  rom[18337] = 16'h83a8;
  rom[18338] = 16'hc50b;
  rom[18339] = 16'he54a;
  rom[18340] = 16'hfd6a;
  rom[18341] = 16'hfce8;
  rom[18342] = 16'hfd49;
  rom[18343] = 16'hf527;
  rom[18344] = 16'hfd68;
  rom[18345] = 16'hf527;
  rom[18346] = 16'hf548;
  rom[18347] = 16'hf528;
  rom[18348] = 16'hfd69;
  rom[18349] = 16'hfce8;
  rom[18350] = 16'hecea;
  rom[18351] = 16'habe9;
  rom[18352] = 16'hac8f;
  rom[18353] = 16'hff9e;
  rom[18354] = 16'hffff;
  rom[18355] = 16'hffff;
  rom[18356] = 16'hffff;
  rom[18357] = 16'hffff;
  rom[18358] = 16'hffff;
  rom[18359] = 16'hffff;
  rom[18360] = 16'hffff;
  rom[18361] = 16'hffff;
  rom[18362] = 16'hffff;
  rom[18363] = 16'hffff;
  rom[18364] = 16'hffff;
  rom[18365] = 16'hffff;
  rom[18366] = 16'hffff;
  rom[18367] = 16'hffff;
  rom[18368] = 16'hffff;
  rom[18369] = 16'hffff;
  rom[18370] = 16'hffff;
  rom[18371] = 16'hffff;
  rom[18372] = 16'hffff;
  rom[18373] = 16'hffff;
  rom[18374] = 16'hffff;
  rom[18375] = 16'hffff;
  rom[18376] = 16'hffff;
  rom[18377] = 16'hffff;
  rom[18378] = 16'hffff;
  rom[18379] = 16'hffff;
  rom[18380] = 16'hffff;
  rom[18381] = 16'hffff;
  rom[18382] = 16'hffff;
  rom[18383] = 16'hffff;
  rom[18384] = 16'hffff;
  rom[18385] = 16'hffff;
  rom[18386] = 16'hffff;
  rom[18387] = 16'hffff;
  rom[18388] = 16'hffff;
  rom[18389] = 16'hffff;
  rom[18390] = 16'hffff;
  rom[18391] = 16'hffff;
  rom[18392] = 16'hffff;
  rom[18393] = 16'hffff;
  rom[18394] = 16'hffff;
  rom[18395] = 16'hffff;
  rom[18396] = 16'hffff;
  rom[18397] = 16'hffff;
  rom[18398] = 16'hffff;
  rom[18399] = 16'hffff;
  rom[18400] = 16'hffff;
  rom[18401] = 16'hffff;
  rom[18402] = 16'hffff;
  rom[18403] = 16'hffff;
  rom[18404] = 16'hffff;
  rom[18405] = 16'hffff;
  rom[18406] = 16'hffff;
  rom[18407] = 16'hffff;
  rom[18408] = 16'hffff;
  rom[18409] = 16'hffff;
  rom[18410] = 16'hffff;
  rom[18411] = 16'hffff;
  rom[18412] = 16'hffff;
  rom[18413] = 16'hffff;
  rom[18414] = 16'hffff;
  rom[18415] = 16'hffff;
  rom[18416] = 16'hffff;
  rom[18417] = 16'hffff;
  rom[18418] = 16'hffff;
  rom[18419] = 16'hffff;
  rom[18420] = 16'hffff;
  rom[18421] = 16'hffff;
  rom[18422] = 16'hffff;
  rom[18423] = 16'hffff;
  rom[18424] = 16'hffff;
  rom[18425] = 16'hffff;
  rom[18426] = 16'he6fa;
  rom[18427] = 16'h5ac3;
  rom[18428] = 16'hd64c;
  rom[18429] = 16'hf70a;
  rom[18430] = 16'hf709;
  rom[18431] = 16'hff4a;
  rom[18432] = 16'hf709;
  rom[18433] = 16'hff29;
  rom[18434] = 16'hff08;
  rom[18435] = 16'hff28;
  rom[18436] = 16'hf708;
  rom[18437] = 16'hff28;
  rom[18438] = 16'hff08;
  rom[18439] = 16'hff28;
  rom[18440] = 16'hf708;
  rom[18441] = 16'hff28;
  rom[18442] = 16'hff08;
  rom[18443] = 16'hff28;
  rom[18444] = 16'hf708;
  rom[18445] = 16'hf729;
  rom[18446] = 16'hf709;
  rom[18447] = 16'hff4c;
  rom[18448] = 16'ha405;
  rom[18449] = 16'h7aa3;
  rom[18450] = 16'hdd6c;
  rom[18451] = 16'hf569;
  rom[18452] = 16'hfd07;
  rom[18453] = 16'hfd09;
  rom[18454] = 16'hf509;
  rom[18455] = 16'hf5ab;
  rom[18456] = 16'hbcaa;
  rom[18457] = 16'h7307;
  rom[18458] = 16'hbd52;
  rom[18459] = 16'hffbe;
  rom[18460] = 16'hffff;
  rom[18461] = 16'hffdf;
  rom[18462] = 16'hffff;
  rom[18463] = 16'hffff;
  rom[18464] = 16'hffdf;
  rom[18465] = 16'hffff;
  rom[18466] = 16'hffff;
  rom[18467] = 16'hffff;
  rom[18468] = 16'hffdf;
  rom[18469] = 16'hffbe;
  rom[18470] = 16'h7bef;
  rom[18471] = 16'h2945;
  rom[18472] = 16'h1061;
  rom[18473] = 16'h18a2;
  rom[18474] = 16'h18a2;
  rom[18475] = 16'h18c3;
  rom[18476] = 16'h18a2;
  rom[18477] = 16'h18a2;
  rom[18478] = 16'h18a2;
  rom[18479] = 16'h18c3;
  rom[18480] = 16'h10c2;
  rom[18481] = 16'h18e3;
  rom[18482] = 16'h10a2;
  rom[18483] = 16'h18c3;
  rom[18484] = 16'h0881;
  rom[18485] = 16'h18c3;
  rom[18486] = 16'h10a2;
  rom[18487] = 16'h9471;
  rom[18488] = 16'hf79e;
  rom[18489] = 16'hffff;
  rom[18490] = 16'hffff;
  rom[18491] = 16'hffff;
  rom[18492] = 16'hffff;
  rom[18493] = 16'hffff;
  rom[18494] = 16'hffff;
  rom[18495] = 16'hffff;
  rom[18496] = 16'hffff;
  rom[18497] = 16'hffff;
  rom[18498] = 16'hffff;
  rom[18499] = 16'hffff;
  rom[18500] = 16'hffff;
  rom[18501] = 16'hffff;
  rom[18502] = 16'hffff;
  rom[18503] = 16'hffff;
  rom[18504] = 16'hffff;
  rom[18505] = 16'hffdf;
  rom[18506] = 16'hce39;
  rom[18507] = 16'h5aaa;
  rom[18508] = 16'h0881;
  rom[18509] = 16'h10a2;
  rom[18510] = 16'h1082;
  rom[18511] = 16'h18a2;
  rom[18512] = 16'h10a2;
  rom[18513] = 16'h18c3;
  rom[18514] = 16'h18a2;
  rom[18515] = 16'h20c3;
  rom[18516] = 16'h1061;
  rom[18517] = 16'h18c3;
  rom[18518] = 16'h18a2;
  rom[18519] = 16'h18a3;
  rom[18520] = 16'h18a2;
  rom[18521] = 16'h18a2;
  rom[18522] = 16'h10a2;
  rom[18523] = 16'h4a49;
  rom[18524] = 16'hbdb6;
  rom[18525] = 16'hffff;
  rom[18526] = 16'hffff;
  rom[18527] = 16'hffff;
  rom[18528] = 16'hffff;
  rom[18529] = 16'hffff;
  rom[18530] = 16'hffff;
  rom[18531] = 16'hffdf;
  rom[18532] = 16'hffff;
  rom[18533] = 16'hffff;
  rom[18534] = 16'hffff;
  rom[18535] = 16'heefa;
  rom[18536] = 16'h8bab;
  rom[18537] = 16'ha409;
  rom[18538] = 16'hdd8c;
  rom[18539] = 16'hf549;
  rom[18540] = 16'hfd08;
  rom[18541] = 16'hfd49;
  rom[18542] = 16'hfd28;
  rom[18543] = 16'hf547;
  rom[18544] = 16'hed47;
  rom[18545] = 16'hf548;
  rom[18546] = 16'hf529;
  rom[18547] = 16'hf529;
  rom[18548] = 16'hf4e8;
  rom[18549] = 16'hfd4a;
  rom[18550] = 16'he52c;
  rom[18551] = 16'h9368;
  rom[18552] = 16'hcdd5;
  rom[18553] = 16'hffff;
  rom[18554] = 16'hffff;
  rom[18555] = 16'hffff;
  rom[18556] = 16'hffff;
  rom[18557] = 16'hffff;
  rom[18558] = 16'hffff;
  rom[18559] = 16'hffff;
  rom[18560] = 16'hffff;
  rom[18561] = 16'hffff;
  rom[18562] = 16'hffff;
  rom[18563] = 16'hffff;
  rom[18564] = 16'hffff;
  rom[18565] = 16'hffff;
  rom[18566] = 16'hffff;
  rom[18567] = 16'hffff;
  rom[18568] = 16'hffff;
  rom[18569] = 16'hffff;
  rom[18570] = 16'hffff;
  rom[18571] = 16'hffff;
  rom[18572] = 16'hffff;
  rom[18573] = 16'hffff;
  rom[18574] = 16'hffff;
  rom[18575] = 16'hffff;
  rom[18576] = 16'hffff;
  rom[18577] = 16'hffff;
  rom[18578] = 16'hffff;
  rom[18579] = 16'hffff;
  rom[18580] = 16'hffff;
  rom[18581] = 16'hffff;
  rom[18582] = 16'hffff;
  rom[18583] = 16'hffff;
  rom[18584] = 16'hffff;
  rom[18585] = 16'hffff;
  rom[18586] = 16'hffff;
  rom[18587] = 16'hffff;
  rom[18588] = 16'hffff;
  rom[18589] = 16'hffff;
  rom[18590] = 16'hffff;
  rom[18591] = 16'hffff;
  rom[18592] = 16'hffff;
  rom[18593] = 16'hffff;
  rom[18594] = 16'hffff;
  rom[18595] = 16'hffff;
  rom[18596] = 16'hffff;
  rom[18597] = 16'hffff;
  rom[18598] = 16'hffff;
  rom[18599] = 16'hffff;
  rom[18600] = 16'hffff;
  rom[18601] = 16'hffff;
  rom[18602] = 16'hffff;
  rom[18603] = 16'hffff;
  rom[18604] = 16'hffff;
  rom[18605] = 16'hffff;
  rom[18606] = 16'hffff;
  rom[18607] = 16'hffff;
  rom[18608] = 16'hffff;
  rom[18609] = 16'hffff;
  rom[18610] = 16'hffff;
  rom[18611] = 16'hffff;
  rom[18612] = 16'hffff;
  rom[18613] = 16'hffff;
  rom[18614] = 16'hffff;
  rom[18615] = 16'hffff;
  rom[18616] = 16'hffff;
  rom[18617] = 16'hffff;
  rom[18618] = 16'hffff;
  rom[18619] = 16'hffff;
  rom[18620] = 16'hffff;
  rom[18621] = 16'hffff;
  rom[18622] = 16'hffff;
  rom[18623] = 16'hffff;
  rom[18624] = 16'hffff;
  rom[18625] = 16'hffdf;
  rom[18626] = 16'hffbe;
  rom[18627] = 16'h5ac5;
  rom[18628] = 16'hcdec;
  rom[18629] = 16'hf72c;
  rom[18630] = 16'hff4a;
  rom[18631] = 16'hff29;
  rom[18632] = 16'hf72a;
  rom[18633] = 16'hf729;
  rom[18634] = 16'hff29;
  rom[18635] = 16'hff28;
  rom[18636] = 16'hff29;
  rom[18637] = 16'hff28;
  rom[18638] = 16'hff29;
  rom[18639] = 16'hff28;
  rom[18640] = 16'hff29;
  rom[18641] = 16'hff28;
  rom[18642] = 16'hff29;
  rom[18643] = 16'hff28;
  rom[18644] = 16'hff2a;
  rom[18645] = 16'hf729;
  rom[18646] = 16'hff4b;
  rom[18647] = 16'hfeea;
  rom[18648] = 16'hf68d;
  rom[18649] = 16'h6a61;
  rom[18650] = 16'hccca;
  rom[18651] = 16'he549;
  rom[18652] = 16'hfd49;
  rom[18653] = 16'hfd28;
  rom[18654] = 16'hfd08;
  rom[18655] = 16'hf568;
  rom[18656] = 16'hed6c;
  rom[18657] = 16'hbcab;
  rom[18658] = 16'h7b07;
  rom[18659] = 16'hcdf5;
  rom[18660] = 16'hffff;
  rom[18661] = 16'hffff;
  rom[18662] = 16'hffff;
  rom[18663] = 16'hffff;
  rom[18664] = 16'hffff;
  rom[18665] = 16'hffff;
  rom[18666] = 16'hffff;
  rom[18667] = 16'hffff;
  rom[18668] = 16'hffff;
  rom[18669] = 16'hffbe;
  rom[18670] = 16'hff9e;
  rom[18671] = 16'h8c31;
  rom[18672] = 16'h20e4;
  rom[18673] = 16'h20e3;
  rom[18674] = 16'h20e3;
  rom[18675] = 16'h1882;
  rom[18676] = 16'h20e3;
  rom[18677] = 16'h20e3;
  rom[18678] = 16'h18a2;
  rom[18679] = 16'h18c3;
  rom[18680] = 16'h20e3;
  rom[18681] = 16'h0840;
  rom[18682] = 16'h1082;
  rom[18683] = 16'h18c2;
  rom[18684] = 16'h2124;
  rom[18685] = 16'h2103;
  rom[18686] = 16'had34;
  rom[18687] = 16'hef3c;
  rom[18688] = 16'hffff;
  rom[18689] = 16'hffff;
  rom[18690] = 16'hffff;
  rom[18691] = 16'hffff;
  rom[18692] = 16'hffff;
  rom[18693] = 16'hffff;
  rom[18694] = 16'hffff;
  rom[18695] = 16'hffff;
  rom[18696] = 16'hffff;
  rom[18697] = 16'hffff;
  rom[18698] = 16'hffff;
  rom[18699] = 16'hffff;
  rom[18700] = 16'hffff;
  rom[18701] = 16'hffff;
  rom[18702] = 16'hffff;
  rom[18703] = 16'hffff;
  rom[18704] = 16'hffff;
  rom[18705] = 16'hffff;
  rom[18706] = 16'hffff;
  rom[18707] = 16'hc5f8;
  rom[18708] = 16'h5acb;
  rom[18709] = 16'h20e3;
  rom[18710] = 16'h2103;
  rom[18711] = 16'h10a2;
  rom[18712] = 16'h1081;
  rom[18713] = 16'h18a2;
  rom[18714] = 16'h1062;
  rom[18715] = 16'h20c3;
  rom[18716] = 16'h2924;
  rom[18717] = 16'h18c3;
  rom[18718] = 16'h20c3;
  rom[18719] = 16'h20e3;
  rom[18720] = 16'h18a2;
  rom[18721] = 16'h18c3;
  rom[18722] = 16'h5249;
  rom[18723] = 16'hce39;
  rom[18724] = 16'hffff;
  rom[18725] = 16'hffdf;
  rom[18726] = 16'hffff;
  rom[18727] = 16'hffff;
  rom[18728] = 16'hffff;
  rom[18729] = 16'hffff;
  rom[18730] = 16'hffff;
  rom[18731] = 16'hffff;
  rom[18732] = 16'hffdf;
  rom[18733] = 16'hffff;
  rom[18734] = 16'hff7b;
  rom[18735] = 16'ha44d;
  rom[18736] = 16'h82e5;
  rom[18737] = 16'hc4ca;
  rom[18738] = 16'hf58b;
  rom[18739] = 16'hfd69;
  rom[18740] = 16'hfd28;
  rom[18741] = 16'hfd48;
  rom[18742] = 16'hfd48;
  rom[18743] = 16'hf527;
  rom[18744] = 16'hf548;
  rom[18745] = 16'hf528;
  rom[18746] = 16'hfd49;
  rom[18747] = 16'hfd29;
  rom[18748] = 16'hfd4a;
  rom[18749] = 16'he50a;
  rom[18750] = 16'hc44b;
  rom[18751] = 16'h93aa;
  rom[18752] = 16'hef1a;
  rom[18753] = 16'hffff;
  rom[18754] = 16'hffff;
  rom[18755] = 16'hffff;
  rom[18756] = 16'hffff;
  rom[18757] = 16'hffff;
  rom[18758] = 16'hffff;
  rom[18759] = 16'hffff;
  rom[18760] = 16'hffff;
  rom[18761] = 16'hffff;
  rom[18762] = 16'hffff;
  rom[18763] = 16'hffff;
  rom[18764] = 16'hffff;
  rom[18765] = 16'hffff;
  rom[18766] = 16'hffff;
  rom[18767] = 16'hffff;
  rom[18768] = 16'hffff;
  rom[18769] = 16'hffff;
  rom[18770] = 16'hffff;
  rom[18771] = 16'hffff;
  rom[18772] = 16'hffff;
  rom[18773] = 16'hffff;
  rom[18774] = 16'hffff;
  rom[18775] = 16'hffff;
  rom[18776] = 16'hffff;
  rom[18777] = 16'hffff;
  rom[18778] = 16'hffff;
  rom[18779] = 16'hffff;
  rom[18780] = 16'hffff;
  rom[18781] = 16'hffff;
  rom[18782] = 16'hffff;
  rom[18783] = 16'hffff;
  rom[18784] = 16'hffff;
  rom[18785] = 16'hffff;
  rom[18786] = 16'hffff;
  rom[18787] = 16'hffff;
  rom[18788] = 16'hffff;
  rom[18789] = 16'hffff;
  rom[18790] = 16'hffff;
  rom[18791] = 16'hffff;
  rom[18792] = 16'hffff;
  rom[18793] = 16'hffff;
  rom[18794] = 16'hffff;
  rom[18795] = 16'hffff;
  rom[18796] = 16'hffff;
  rom[18797] = 16'hffff;
  rom[18798] = 16'hffff;
  rom[18799] = 16'hffff;
  rom[18800] = 16'hffff;
  rom[18801] = 16'hffff;
  rom[18802] = 16'hffff;
  rom[18803] = 16'hffff;
  rom[18804] = 16'hffff;
  rom[18805] = 16'hffff;
  rom[18806] = 16'hffff;
  rom[18807] = 16'hffff;
  rom[18808] = 16'hffff;
  rom[18809] = 16'hffff;
  rom[18810] = 16'hffff;
  rom[18811] = 16'hffff;
  rom[18812] = 16'hffff;
  rom[18813] = 16'hffff;
  rom[18814] = 16'hffff;
  rom[18815] = 16'hffff;
  rom[18816] = 16'hffff;
  rom[18817] = 16'hffff;
  rom[18818] = 16'hffff;
  rom[18819] = 16'hffff;
  rom[18820] = 16'hffff;
  rom[18821] = 16'hffff;
  rom[18822] = 16'hffff;
  rom[18823] = 16'hffff;
  rom[18824] = 16'hffdf;
  rom[18825] = 16'hffff;
  rom[18826] = 16'hf77d;
  rom[18827] = 16'h6b28;
  rom[18828] = 16'hc5ed;
  rom[18829] = 16'hff4d;
  rom[18830] = 16'hef28;
  rom[18831] = 16'hf749;
  rom[18832] = 16'hf728;
  rom[18833] = 16'hf729;
  rom[18834] = 16'hf728;
  rom[18835] = 16'hff28;
  rom[18836] = 16'hff08;
  rom[18837] = 16'hff28;
  rom[18838] = 16'hf708;
  rom[18839] = 16'hff28;
  rom[18840] = 16'hff08;
  rom[18841] = 16'hff28;
  rom[18842] = 16'hf708;
  rom[18843] = 16'hff28;
  rom[18844] = 16'hff09;
  rom[18845] = 16'hff29;
  rom[18846] = 16'hf709;
  rom[18847] = 16'hf6ea;
  rom[18848] = 16'hf6ec;
  rom[18849] = 16'h93a5;
  rom[18850] = 16'h6a61;
  rom[18851] = 16'he54a;
  rom[18852] = 16'hf529;
  rom[18853] = 16'hfd28;
  rom[18854] = 16'hfd27;
  rom[18855] = 16'hfd48;
  rom[18856] = 16'hed49;
  rom[18857] = 16'he58d;
  rom[18858] = 16'hb46a;
  rom[18859] = 16'h7ae6;
  rom[18860] = 16'hc5b3;
  rom[18861] = 16'hff9d;
  rom[18862] = 16'hffdf;
  rom[18863] = 16'hffff;
  rom[18864] = 16'hffdf;
  rom[18865] = 16'hffff;
  rom[18866] = 16'hffff;
  rom[18867] = 16'hffff;
  rom[18868] = 16'hffff;
  rom[18869] = 16'hffff;
  rom[18870] = 16'hffdf;
  rom[18871] = 16'hffbf;
  rom[18872] = 16'hbd96;
  rom[18873] = 16'h62cb;
  rom[18874] = 16'h18c2;
  rom[18875] = 16'h18a2;
  rom[18876] = 16'h1082;
  rom[18877] = 16'h20c3;
  rom[18878] = 16'h1082;
  rom[18879] = 16'h18c3;
  rom[18880] = 16'h10a2;
  rom[18881] = 16'h2104;
  rom[18882] = 16'h18c3;
  rom[18883] = 16'h2104;
  rom[18884] = 16'h5269;
  rom[18885] = 16'hbdb7;
  rom[18886] = 16'hf7be;
  rom[18887] = 16'hffff;
  rom[18888] = 16'hffff;
  rom[18889] = 16'hffff;
  rom[18890] = 16'hffff;
  rom[18891] = 16'hffff;
  rom[18892] = 16'hffff;
  rom[18893] = 16'hffff;
  rom[18894] = 16'hffff;
  rom[18895] = 16'hffff;
  rom[18896] = 16'hffff;
  rom[18897] = 16'hffff;
  rom[18898] = 16'hffff;
  rom[18899] = 16'hffff;
  rom[18900] = 16'hffff;
  rom[18901] = 16'hffff;
  rom[18902] = 16'hffff;
  rom[18903] = 16'hffdf;
  rom[18904] = 16'hffff;
  rom[18905] = 16'hffdf;
  rom[18906] = 16'hffff;
  rom[18907] = 16'hffff;
  rom[18908] = 16'hdebb;
  rom[18909] = 16'h9471;
  rom[18910] = 16'h3186;
  rom[18911] = 16'h18e3;
  rom[18912] = 16'h10a2;
  rom[18913] = 16'h18a3;
  rom[18914] = 16'h18c3;
  rom[18915] = 16'h10a2;
  rom[18916] = 16'h1082;
  rom[18917] = 16'h18c3;
  rom[18918] = 16'h18a2;
  rom[18919] = 16'h18a3;
  rom[18920] = 16'h3986;
  rom[18921] = 16'h8c30;
  rom[18922] = 16'he6fb;
  rom[18923] = 16'hffdf;
  rom[18924] = 16'hffbf;
  rom[18925] = 16'hffff;
  rom[18926] = 16'hffdf;
  rom[18927] = 16'hffff;
  rom[18928] = 16'hffdf;
  rom[18929] = 16'hffff;
  rom[18930] = 16'hffdf;
  rom[18931] = 16'hffff;
  rom[18932] = 16'hffbe;
  rom[18933] = 16'hff9c;
  rom[18934] = 16'h93cb;
  rom[18935] = 16'h8b26;
  rom[18936] = 16'hd52b;
  rom[18937] = 16'hed8b;
  rom[18938] = 16'hf548;
  rom[18939] = 16'hfd07;
  rom[18940] = 16'hfd07;
  rom[18941] = 16'hfd07;
  rom[18942] = 16'hf527;
  rom[18943] = 16'hf547;
  rom[18944] = 16'hf548;
  rom[18945] = 16'hfd28;
  rom[18946] = 16'hfd08;
  rom[18947] = 16'hfd08;
  rom[18948] = 16'hed2a;
  rom[18949] = 16'he54c;
  rom[18950] = 16'h82e5;
  rom[18951] = 16'hb4f1;
  rom[18952] = 16'hffbd;
  rom[18953] = 16'hffff;
  rom[18954] = 16'hffff;
  rom[18955] = 16'hffff;
  rom[18956] = 16'hffff;
  rom[18957] = 16'hffff;
  rom[18958] = 16'hffff;
  rom[18959] = 16'hffff;
  rom[18960] = 16'hffff;
  rom[18961] = 16'hffff;
  rom[18962] = 16'hffff;
  rom[18963] = 16'hffff;
  rom[18964] = 16'hffff;
  rom[18965] = 16'hffff;
  rom[18966] = 16'hffff;
  rom[18967] = 16'hffff;
  rom[18968] = 16'hffff;
  rom[18969] = 16'hffff;
  rom[18970] = 16'hffff;
  rom[18971] = 16'hffff;
  rom[18972] = 16'hffff;
  rom[18973] = 16'hffff;
  rom[18974] = 16'hffff;
  rom[18975] = 16'hffff;
  rom[18976] = 16'hffff;
  rom[18977] = 16'hffff;
  rom[18978] = 16'hffff;
  rom[18979] = 16'hffff;
  rom[18980] = 16'hffff;
  rom[18981] = 16'hffff;
  rom[18982] = 16'hffff;
  rom[18983] = 16'hffff;
  rom[18984] = 16'hffff;
  rom[18985] = 16'hffff;
  rom[18986] = 16'hffff;
  rom[18987] = 16'hffff;
  rom[18988] = 16'hffff;
  rom[18989] = 16'hffff;
  rom[18990] = 16'hffff;
  rom[18991] = 16'hffff;
  rom[18992] = 16'hffff;
  rom[18993] = 16'hffff;
  rom[18994] = 16'hffff;
  rom[18995] = 16'hffff;
  rom[18996] = 16'hffff;
  rom[18997] = 16'hffff;
  rom[18998] = 16'hffff;
  rom[18999] = 16'hffff;
  rom[19000] = 16'hffff;
  rom[19001] = 16'hffff;
  rom[19002] = 16'hffff;
  rom[19003] = 16'hffff;
  rom[19004] = 16'hffff;
  rom[19005] = 16'hffff;
  rom[19006] = 16'hffff;
  rom[19007] = 16'hffff;
  rom[19008] = 16'hffff;
  rom[19009] = 16'hffff;
  rom[19010] = 16'hffff;
  rom[19011] = 16'hffff;
  rom[19012] = 16'hffff;
  rom[19013] = 16'hffff;
  rom[19014] = 16'hffff;
  rom[19015] = 16'hffff;
  rom[19016] = 16'hffff;
  rom[19017] = 16'hffff;
  rom[19018] = 16'hffff;
  rom[19019] = 16'hffff;
  rom[19020] = 16'hffff;
  rom[19021] = 16'hffff;
  rom[19022] = 16'hffff;
  rom[19023] = 16'hffff;
  rom[19024] = 16'hffff;
  rom[19025] = 16'hffff;
  rom[19026] = 16'hffdf;
  rom[19027] = 16'h946e;
  rom[19028] = 16'haccb;
  rom[19029] = 16'he6cb;
  rom[19030] = 16'hff49;
  rom[19031] = 16'hf727;
  rom[19032] = 16'hff49;
  rom[19033] = 16'hff48;
  rom[19034] = 16'hff29;
  rom[19035] = 16'hff28;
  rom[19036] = 16'hff29;
  rom[19037] = 16'hff28;
  rom[19038] = 16'hff29;
  rom[19039] = 16'hff28;
  rom[19040] = 16'hff29;
  rom[19041] = 16'hff28;
  rom[19042] = 16'hff29;
  rom[19043] = 16'hff28;
  rom[19044] = 16'hff2a;
  rom[19045] = 16'hff28;
  rom[19046] = 16'hff0a;
  rom[19047] = 16'hff2b;
  rom[19048] = 16'hf6cb;
  rom[19049] = 16'hd5ea;
  rom[19050] = 16'h5180;
  rom[19051] = 16'hc469;
  rom[19052] = 16'hf54c;
  rom[19053] = 16'hf508;
  rom[19054] = 16'hfd06;
  rom[19055] = 16'hfd89;
  rom[19056] = 16'hfd28;
  rom[19057] = 16'hed29;
  rom[19058] = 16'hed8c;
  rom[19059] = 16'hbc6a;
  rom[19060] = 16'h7264;
  rom[19061] = 16'hc593;
  rom[19062] = 16'hffff;
  rom[19063] = 16'hffff;
  rom[19064] = 16'hffff;
  rom[19065] = 16'hffff;
  rom[19066] = 16'hffff;
  rom[19067] = 16'hffff;
  rom[19068] = 16'hffff;
  rom[19069] = 16'hffff;
  rom[19070] = 16'hffff;
  rom[19071] = 16'hffff;
  rom[19072] = 16'hffdf;
  rom[19073] = 16'hef3d;
  rom[19074] = 16'hce18;
  rom[19075] = 16'h6b4d;
  rom[19076] = 16'h2925;
  rom[19077] = 16'h1082;
  rom[19078] = 16'h1082;
  rom[19079] = 16'h18a3;
  rom[19080] = 16'h18c3;
  rom[19081] = 16'h18c3;
  rom[19082] = 16'h6b0c;
  rom[19083] = 16'hbdf7;
  rom[19084] = 16'hffbf;
  rom[19085] = 16'hffdf;
  rom[19086] = 16'hffff;
  rom[19087] = 16'hffdf;
  rom[19088] = 16'hffff;
  rom[19089] = 16'hffff;
  rom[19090] = 16'hffff;
  rom[19091] = 16'hffff;
  rom[19092] = 16'hffff;
  rom[19093] = 16'hffff;
  rom[19094] = 16'hffff;
  rom[19095] = 16'hffff;
  rom[19096] = 16'hffff;
  rom[19097] = 16'hffff;
  rom[19098] = 16'hffff;
  rom[19099] = 16'hffff;
  rom[19100] = 16'hffff;
  rom[19101] = 16'hffff;
  rom[19102] = 16'hffff;
  rom[19103] = 16'hffff;
  rom[19104] = 16'hffff;
  rom[19105] = 16'hffff;
  rom[19106] = 16'hffff;
  rom[19107] = 16'hffff;
  rom[19108] = 16'hffff;
  rom[19109] = 16'hff9f;
  rom[19110] = 16'hef5d;
  rom[19111] = 16'ha514;
  rom[19112] = 16'h4208;
  rom[19113] = 16'h20e3;
  rom[19114] = 16'h18a3;
  rom[19115] = 16'h18c2;
  rom[19116] = 16'h20e4;
  rom[19117] = 16'h1082;
  rom[19118] = 16'h4208;
  rom[19119] = 16'h9cb3;
  rom[19120] = 16'hef1d;
  rom[19121] = 16'hff9f;
  rom[19122] = 16'hffff;
  rom[19123] = 16'hffdf;
  rom[19124] = 16'hffff;
  rom[19125] = 16'hffbf;
  rom[19126] = 16'hffff;
  rom[19127] = 16'hffdf;
  rom[19128] = 16'hffdf;
  rom[19129] = 16'hffff;
  rom[19130] = 16'hffff;
  rom[19131] = 16'hffde;
  rom[19132] = 16'hf73b;
  rom[19133] = 16'h6a65;
  rom[19134] = 16'h9b88;
  rom[19135] = 16'hd50b;
  rom[19136] = 16'hf58b;
  rom[19137] = 16'hf548;
  rom[19138] = 16'hfd28;
  rom[19139] = 16'hfd27;
  rom[19140] = 16'hfd08;
  rom[19141] = 16'hfd28;
  rom[19142] = 16'hfd68;
  rom[19143] = 16'hf527;
  rom[19144] = 16'hfd48;
  rom[19145] = 16'hfce8;
  rom[19146] = 16'hfd09;
  rom[19147] = 16'hfd08;
  rom[19148] = 16'hf54c;
  rom[19149] = 16'hc46a;
  rom[19150] = 16'h72a6;
  rom[19151] = 16'hde98;
  rom[19152] = 16'hffff;
  rom[19153] = 16'hffff;
  rom[19154] = 16'hffff;
  rom[19155] = 16'hffff;
  rom[19156] = 16'hffff;
  rom[19157] = 16'hffff;
  rom[19158] = 16'hffff;
  rom[19159] = 16'hffff;
  rom[19160] = 16'hffff;
  rom[19161] = 16'hffff;
  rom[19162] = 16'hffff;
  rom[19163] = 16'hffff;
  rom[19164] = 16'hffff;
  rom[19165] = 16'hffff;
  rom[19166] = 16'hffff;
  rom[19167] = 16'hffff;
  rom[19168] = 16'hffff;
  rom[19169] = 16'hffff;
  rom[19170] = 16'hffff;
  rom[19171] = 16'hffff;
  rom[19172] = 16'hffff;
  rom[19173] = 16'hffff;
  rom[19174] = 16'hffff;
  rom[19175] = 16'hffff;
  rom[19176] = 16'hffff;
  rom[19177] = 16'hffff;
  rom[19178] = 16'hffff;
  rom[19179] = 16'hffff;
  rom[19180] = 16'hffff;
  rom[19181] = 16'hffff;
  rom[19182] = 16'hffff;
  rom[19183] = 16'hffff;
  rom[19184] = 16'hffff;
  rom[19185] = 16'hffff;
  rom[19186] = 16'hffff;
  rom[19187] = 16'hffff;
  rom[19188] = 16'hffff;
  rom[19189] = 16'hffff;
  rom[19190] = 16'hffff;
  rom[19191] = 16'hffff;
  rom[19192] = 16'hffff;
  rom[19193] = 16'hffff;
  rom[19194] = 16'hffff;
  rom[19195] = 16'hffff;
  rom[19196] = 16'hffff;
  rom[19197] = 16'hffff;
  rom[19198] = 16'hffff;
  rom[19199] = 16'hffff;
  rom[19200] = 16'hffff;
  rom[19201] = 16'hffff;
  rom[19202] = 16'hffff;
  rom[19203] = 16'hffff;
  rom[19204] = 16'hffff;
  rom[19205] = 16'hffff;
  rom[19206] = 16'hffff;
  rom[19207] = 16'hffff;
  rom[19208] = 16'hffff;
  rom[19209] = 16'hffff;
  rom[19210] = 16'hffff;
  rom[19211] = 16'hffff;
  rom[19212] = 16'hffff;
  rom[19213] = 16'hffff;
  rom[19214] = 16'hffff;
  rom[19215] = 16'hffff;
  rom[19216] = 16'hffff;
  rom[19217] = 16'hffff;
  rom[19218] = 16'hffff;
  rom[19219] = 16'hffff;
  rom[19220] = 16'hffff;
  rom[19221] = 16'hffff;
  rom[19222] = 16'hffff;
  rom[19223] = 16'hffff;
  rom[19224] = 16'hfffe;
  rom[19225] = 16'hffff;
  rom[19226] = 16'hffff;
  rom[19227] = 16'hb532;
  rom[19228] = 16'h6b24;
  rom[19229] = 16'hef0e;
  rom[19230] = 16'hf729;
  rom[19231] = 16'hff28;
  rom[19232] = 16'hff08;
  rom[19233] = 16'hf708;
  rom[19234] = 16'hf728;
  rom[19235] = 16'hff49;
  rom[19236] = 16'hf707;
  rom[19237] = 16'hff49;
  rom[19238] = 16'hf728;
  rom[19239] = 16'hff28;
  rom[19240] = 16'hf708;
  rom[19241] = 16'hff28;
  rom[19242] = 16'hff08;
  rom[19243] = 16'hff28;
  rom[19244] = 16'hf708;
  rom[19245] = 16'hff28;
  rom[19246] = 16'hf709;
  rom[19247] = 16'hf70a;
  rom[19248] = 16'hf74c;
  rom[19249] = 16'hf70c;
  rom[19250] = 16'h8362;
  rom[19251] = 16'h82a4;
  rom[19252] = 16'he52c;
  rom[19253] = 16'hf529;
  rom[19254] = 16'hfce6;
  rom[19255] = 16'hfd08;
  rom[19256] = 16'hfd28;
  rom[19257] = 16'hfd89;
  rom[19258] = 16'hf549;
  rom[19259] = 16'hed2b;
  rom[19260] = 16'hd4ed;
  rom[19261] = 16'h7265;
  rom[19262] = 16'h940d;
  rom[19263] = 16'hded9;
  rom[19264] = 16'hf7de;
  rom[19265] = 16'hffff;
  rom[19266] = 16'hffde;
  rom[19267] = 16'hffff;
  rom[19268] = 16'hffdf;
  rom[19269] = 16'hffff;
  rom[19270] = 16'hffff;
  rom[19271] = 16'hffff;
  rom[19272] = 16'hffff;
  rom[19273] = 16'hffff;
  rom[19274] = 16'hffbf;
  rom[19275] = 16'hffff;
  rom[19276] = 16'hffdf;
  rom[19277] = 16'hef3d;
  rom[19278] = 16'hbdb6;
  rom[19279] = 16'hc5f8;
  rom[19280] = 16'hef5d;
  rom[19281] = 16'hffff;
  rom[19282] = 16'hffff;
  rom[19283] = 16'hffff;
  rom[19284] = 16'hffff;
  rom[19285] = 16'hffff;
  rom[19286] = 16'hffff;
  rom[19287] = 16'hffff;
  rom[19288] = 16'hffff;
  rom[19289] = 16'hffff;
  rom[19290] = 16'hffff;
  rom[19291] = 16'hffff;
  rom[19292] = 16'hffff;
  rom[19293] = 16'hffff;
  rom[19294] = 16'hffff;
  rom[19295] = 16'hffff;
  rom[19296] = 16'hffff;
  rom[19297] = 16'hffff;
  rom[19298] = 16'hffff;
  rom[19299] = 16'hffff;
  rom[19300] = 16'hffff;
  rom[19301] = 16'hffff;
  rom[19302] = 16'hffff;
  rom[19303] = 16'hffff;
  rom[19304] = 16'hffff;
  rom[19305] = 16'hffff;
  rom[19306] = 16'hffff;
  rom[19307] = 16'hffff;
  rom[19308] = 16'hffdf;
  rom[19309] = 16'hffff;
  rom[19310] = 16'hffff;
  rom[19311] = 16'hffff;
  rom[19312] = 16'hffdf;
  rom[19313] = 16'hff9f;
  rom[19314] = 16'hd67a;
  rom[19315] = 16'hc5d7;
  rom[19316] = 16'hd69a;
  rom[19317] = 16'hffdf;
  rom[19318] = 16'hffff;
  rom[19319] = 16'hffff;
  rom[19320] = 16'hffff;
  rom[19321] = 16'hffff;
  rom[19322] = 16'hffdf;
  rom[19323] = 16'hffff;
  rom[19324] = 16'hffff;
  rom[19325] = 16'hffff;
  rom[19326] = 16'hffff;
  rom[19327] = 16'hffdf;
  rom[19328] = 16'hffff;
  rom[19329] = 16'hffde;
  rom[19330] = 16'hff7c;
  rom[19331] = 16'hc5b4;
  rom[19332] = 16'h6ac7;
  rom[19333] = 16'hac4a;
  rom[19334] = 16'hdd2b;
  rom[19335] = 16'hed4a;
  rom[19336] = 16'hf528;
  rom[19337] = 16'hfd28;
  rom[19338] = 16'hfd48;
  rom[19339] = 16'hfd29;
  rom[19340] = 16'hf528;
  rom[19341] = 16'hf549;
  rom[19342] = 16'hf528;
  rom[19343] = 16'hfd47;
  rom[19344] = 16'hfd07;
  rom[19345] = 16'hfd07;
  rom[19346] = 16'hfce7;
  rom[19347] = 16'hfd29;
  rom[19348] = 16'hed2b;
  rom[19349] = 16'h9b88;
  rom[19350] = 16'h940d;
  rom[19351] = 16'hffde;
  rom[19352] = 16'hffff;
  rom[19353] = 16'hffff;
  rom[19354] = 16'hffff;
  rom[19355] = 16'hffff;
  rom[19356] = 16'hffff;
  rom[19357] = 16'hffff;
  rom[19358] = 16'hffff;
  rom[19359] = 16'hffff;
  rom[19360] = 16'hffff;
  rom[19361] = 16'hffff;
  rom[19362] = 16'hffff;
  rom[19363] = 16'hffff;
  rom[19364] = 16'hffff;
  rom[19365] = 16'hffff;
  rom[19366] = 16'hffff;
  rom[19367] = 16'hffff;
  rom[19368] = 16'hffff;
  rom[19369] = 16'hffff;
  rom[19370] = 16'hffff;
  rom[19371] = 16'hffff;
  rom[19372] = 16'hffff;
  rom[19373] = 16'hffff;
  rom[19374] = 16'hffff;
  rom[19375] = 16'hffff;
  rom[19376] = 16'hffff;
  rom[19377] = 16'hffff;
  rom[19378] = 16'hffff;
  rom[19379] = 16'hffff;
  rom[19380] = 16'hffff;
  rom[19381] = 16'hffff;
  rom[19382] = 16'hffff;
  rom[19383] = 16'hffff;
  rom[19384] = 16'hffff;
  rom[19385] = 16'hffff;
  rom[19386] = 16'hffff;
  rom[19387] = 16'hffff;
  rom[19388] = 16'hffff;
  rom[19389] = 16'hffff;
  rom[19390] = 16'hffff;
  rom[19391] = 16'hffff;
  rom[19392] = 16'hffff;
  rom[19393] = 16'hffff;
  rom[19394] = 16'hffff;
  rom[19395] = 16'hffff;
  rom[19396] = 16'hffff;
  rom[19397] = 16'hffff;
  rom[19398] = 16'hffff;
  rom[19399] = 16'hffff;
  rom[19400] = 16'hffff;
  rom[19401] = 16'hffff;
  rom[19402] = 16'hffff;
  rom[19403] = 16'hffff;
  rom[19404] = 16'hffff;
  rom[19405] = 16'hffff;
  rom[19406] = 16'hffff;
  rom[19407] = 16'hffff;
  rom[19408] = 16'hffff;
  rom[19409] = 16'hffff;
  rom[19410] = 16'hffff;
  rom[19411] = 16'hffff;
  rom[19412] = 16'hffff;
  rom[19413] = 16'hffff;
  rom[19414] = 16'hffff;
  rom[19415] = 16'hffff;
  rom[19416] = 16'hffff;
  rom[19417] = 16'hffff;
  rom[19418] = 16'hffff;
  rom[19419] = 16'hffff;
  rom[19420] = 16'hffff;
  rom[19421] = 16'hffff;
  rom[19422] = 16'hffff;
  rom[19423] = 16'hffff;
  rom[19424] = 16'hffff;
  rom[19425] = 16'hffff;
  rom[19426] = 16'hffff;
  rom[19427] = 16'hde98;
  rom[19428] = 16'h62a4;
  rom[19429] = 16'hbd8a;
  rom[19430] = 16'hff4d;
  rom[19431] = 16'hff09;
  rom[19432] = 16'hff2a;
  rom[19433] = 16'hf709;
  rom[19434] = 16'hff09;
  rom[19435] = 16'hf708;
  rom[19436] = 16'hff29;
  rom[19437] = 16'hf728;
  rom[19438] = 16'hff49;
  rom[19439] = 16'hff28;
  rom[19440] = 16'hff29;
  rom[19441] = 16'hff28;
  rom[19442] = 16'hff29;
  rom[19443] = 16'hff28;
  rom[19444] = 16'hff29;
  rom[19445] = 16'hff48;
  rom[19446] = 16'hff29;
  rom[19447] = 16'hff0a;
  rom[19448] = 16'heeea;
  rom[19449] = 16'hff4c;
  rom[19450] = 16'he64b;
  rom[19451] = 16'h61e0;
  rom[19452] = 16'hdccc;
  rom[19453] = 16'hed2a;
  rom[19454] = 16'hfd4a;
  rom[19455] = 16'hfd08;
  rom[19456] = 16'hfd28;
  rom[19457] = 16'hfd27;
  rom[19458] = 16'hfd27;
  rom[19459] = 16'hfd4a;
  rom[19460] = 16'hf54c;
  rom[19461] = 16'hd50d;
  rom[19462] = 16'h9bea;
  rom[19463] = 16'h6ac6;
  rom[19464] = 16'ha4d0;
  rom[19465] = 16'hef5a;
  rom[19466] = 16'hffde;
  rom[19467] = 16'hffff;
  rom[19468] = 16'hffff;
  rom[19469] = 16'hffff;
  rom[19470] = 16'hffff;
  rom[19471] = 16'hffff;
  rom[19472] = 16'hffff;
  rom[19473] = 16'hffff;
  rom[19474] = 16'hffff;
  rom[19475] = 16'hffff;
  rom[19476] = 16'hffff;
  rom[19477] = 16'hffff;
  rom[19478] = 16'hffdf;
  rom[19479] = 16'hffff;
  rom[19480] = 16'hffff;
  rom[19481] = 16'hffff;
  rom[19482] = 16'hffff;
  rom[19483] = 16'hffff;
  rom[19484] = 16'hffff;
  rom[19485] = 16'hffff;
  rom[19486] = 16'hffff;
  rom[19487] = 16'hffff;
  rom[19488] = 16'hffff;
  rom[19489] = 16'hffff;
  rom[19490] = 16'hffff;
  rom[19491] = 16'hffff;
  rom[19492] = 16'hffff;
  rom[19493] = 16'hffff;
  rom[19494] = 16'hffff;
  rom[19495] = 16'hffff;
  rom[19496] = 16'hffff;
  rom[19497] = 16'hffff;
  rom[19498] = 16'hffff;
  rom[19499] = 16'hffff;
  rom[19500] = 16'hffdf;
  rom[19501] = 16'hffff;
  rom[19502] = 16'hffff;
  rom[19503] = 16'hffff;
  rom[19504] = 16'hffff;
  rom[19505] = 16'hffff;
  rom[19506] = 16'hffff;
  rom[19507] = 16'hffff;
  rom[19508] = 16'hffff;
  rom[19509] = 16'hffff;
  rom[19510] = 16'hffff;
  rom[19511] = 16'hffff;
  rom[19512] = 16'hffff;
  rom[19513] = 16'hffff;
  rom[19514] = 16'hffff;
  rom[19515] = 16'hffff;
  rom[19516] = 16'hffff;
  rom[19517] = 16'hffff;
  rom[19518] = 16'hffff;
  rom[19519] = 16'hffff;
  rom[19520] = 16'hffff;
  rom[19521] = 16'hffff;
  rom[19522] = 16'hffff;
  rom[19523] = 16'hffff;
  rom[19524] = 16'hffff;
  rom[19525] = 16'hffff;
  rom[19526] = 16'hffff;
  rom[19527] = 16'hffdf;
  rom[19528] = 16'hff7d;
  rom[19529] = 16'hde36;
  rom[19530] = 16'h936a;
  rom[19531] = 16'h82e6;
  rom[19532] = 16'hc4ac;
  rom[19533] = 16'hd52b;
  rom[19534] = 16'hf56b;
  rom[19535] = 16'hf549;
  rom[19536] = 16'hfd07;
  rom[19537] = 16'hfd47;
  rom[19538] = 16'hfd28;
  rom[19539] = 16'hf508;
  rom[19540] = 16'hf56a;
  rom[19541] = 16'hf569;
  rom[19542] = 16'hf528;
  rom[19543] = 16'hfd27;
  rom[19544] = 16'hfd07;
  rom[19545] = 16'hfce7;
  rom[19546] = 16'hfd09;
  rom[19547] = 16'hf52a;
  rom[19548] = 16'hcc6a;
  rom[19549] = 16'h8b48;
  rom[19550] = 16'hf77b;
  rom[19551] = 16'hfffe;
  rom[19552] = 16'hffff;
  rom[19553] = 16'hffff;
  rom[19554] = 16'hffff;
  rom[19555] = 16'hffff;
  rom[19556] = 16'hffff;
  rom[19557] = 16'hffff;
  rom[19558] = 16'hffff;
  rom[19559] = 16'hffff;
  rom[19560] = 16'hffff;
  rom[19561] = 16'hffff;
  rom[19562] = 16'hffff;
  rom[19563] = 16'hffff;
  rom[19564] = 16'hffff;
  rom[19565] = 16'hffff;
  rom[19566] = 16'hffff;
  rom[19567] = 16'hffff;
  rom[19568] = 16'hffff;
  rom[19569] = 16'hffff;
  rom[19570] = 16'hffff;
  rom[19571] = 16'hffff;
  rom[19572] = 16'hffff;
  rom[19573] = 16'hffff;
  rom[19574] = 16'hffff;
  rom[19575] = 16'hffff;
  rom[19576] = 16'hffff;
  rom[19577] = 16'hffff;
  rom[19578] = 16'hffff;
  rom[19579] = 16'hffff;
  rom[19580] = 16'hffff;
  rom[19581] = 16'hffff;
  rom[19582] = 16'hffff;
  rom[19583] = 16'hffff;
  rom[19584] = 16'hffff;
  rom[19585] = 16'hffff;
  rom[19586] = 16'hffff;
  rom[19587] = 16'hffff;
  rom[19588] = 16'hffff;
  rom[19589] = 16'hffff;
  rom[19590] = 16'hffff;
  rom[19591] = 16'hffff;
  rom[19592] = 16'hffff;
  rom[19593] = 16'hffff;
  rom[19594] = 16'hffff;
  rom[19595] = 16'hffff;
  rom[19596] = 16'hffff;
  rom[19597] = 16'hffff;
  rom[19598] = 16'hffff;
  rom[19599] = 16'hffff;
  rom[19600] = 16'hffff;
  rom[19601] = 16'hffff;
  rom[19602] = 16'hffff;
  rom[19603] = 16'hffff;
  rom[19604] = 16'hffff;
  rom[19605] = 16'hffff;
  rom[19606] = 16'hffff;
  rom[19607] = 16'hffff;
  rom[19608] = 16'hffff;
  rom[19609] = 16'hffff;
  rom[19610] = 16'hffff;
  rom[19611] = 16'hffff;
  rom[19612] = 16'hffff;
  rom[19613] = 16'hffff;
  rom[19614] = 16'hffff;
  rom[19615] = 16'hffff;
  rom[19616] = 16'hffff;
  rom[19617] = 16'hffff;
  rom[19618] = 16'hffff;
  rom[19619] = 16'hffff;
  rom[19620] = 16'hffff;
  rom[19621] = 16'hffff;
  rom[19622] = 16'hffff;
  rom[19623] = 16'hffff;
  rom[19624] = 16'hffff;
  rom[19625] = 16'hffff;
  rom[19626] = 16'hffdf;
  rom[19627] = 16'hff9d;
  rom[19628] = 16'h8beb;
  rom[19629] = 16'h7344;
  rom[19630] = 16'hce2b;
  rom[19631] = 16'hff2d;
  rom[19632] = 16'hf6eb;
  rom[19633] = 16'hff0b;
  rom[19634] = 16'hf76a;
  rom[19635] = 16'hf728;
  rom[19636] = 16'hff49;
  rom[19637] = 16'hf709;
  rom[19638] = 16'hf708;
  rom[19639] = 16'hff28;
  rom[19640] = 16'hff08;
  rom[19641] = 16'hff28;
  rom[19642] = 16'hf708;
  rom[19643] = 16'hff28;
  rom[19644] = 16'hff08;
  rom[19645] = 16'hff28;
  rom[19646] = 16'hf728;
  rom[19647] = 16'hff4b;
  rom[19648] = 16'heec9;
  rom[19649] = 16'hff4b;
  rom[19650] = 16'hf6eb;
  rom[19651] = 16'h9386;
  rom[19652] = 16'h8aa3;
  rom[19653] = 16'he50b;
  rom[19654] = 16'hece8;
  rom[19655] = 16'hfd29;
  rom[19656] = 16'hfd27;
  rom[19657] = 16'hfd47;
  rom[19658] = 16'hfd47;
  rom[19659] = 16'hfd28;
  rom[19660] = 16'hf529;
  rom[19661] = 16'hf54c;
  rom[19662] = 16'he54d;
  rom[19663] = 16'hcd2d;
  rom[19664] = 16'h6ac4;
  rom[19665] = 16'h6ae7;
  rom[19666] = 16'ha4d1;
  rom[19667] = 16'hffff;
  rom[19668] = 16'hffff;
  rom[19669] = 16'hffff;
  rom[19670] = 16'hffff;
  rom[19671] = 16'hffff;
  rom[19672] = 16'hffff;
  rom[19673] = 16'hffff;
  rom[19674] = 16'hffff;
  rom[19675] = 16'hffff;
  rom[19676] = 16'hffff;
  rom[19677] = 16'hffff;
  rom[19678] = 16'hffff;
  rom[19679] = 16'hffff;
  rom[19680] = 16'hffff;
  rom[19681] = 16'hffff;
  rom[19682] = 16'hffff;
  rom[19683] = 16'hffff;
  rom[19684] = 16'hffff;
  rom[19685] = 16'hffff;
  rom[19686] = 16'hffff;
  rom[19687] = 16'hffff;
  rom[19688] = 16'hffff;
  rom[19689] = 16'hffff;
  rom[19690] = 16'hffff;
  rom[19691] = 16'hffff;
  rom[19692] = 16'hffff;
  rom[19693] = 16'hffff;
  rom[19694] = 16'hffdf;
  rom[19695] = 16'hff9e;
  rom[19696] = 16'hd69a;
  rom[19697] = 16'hd65a;
  rom[19698] = 16'hf79e;
  rom[19699] = 16'hffdf;
  rom[19700] = 16'hffff;
  rom[19701] = 16'hffff;
  rom[19702] = 16'hffff;
  rom[19703] = 16'hffff;
  rom[19704] = 16'hffff;
  rom[19705] = 16'hffff;
  rom[19706] = 16'hffff;
  rom[19707] = 16'hffff;
  rom[19708] = 16'hffff;
  rom[19709] = 16'hffff;
  rom[19710] = 16'hffff;
  rom[19711] = 16'hffff;
  rom[19712] = 16'hffff;
  rom[19713] = 16'hffff;
  rom[19714] = 16'hffff;
  rom[19715] = 16'hffff;
  rom[19716] = 16'hffff;
  rom[19717] = 16'hffff;
  rom[19718] = 16'hffff;
  rom[19719] = 16'hffff;
  rom[19720] = 16'hffff;
  rom[19721] = 16'hffff;
  rom[19722] = 16'hffff;
  rom[19723] = 16'hffff;
  rom[19724] = 16'hffff;
  rom[19725] = 16'hffff;
  rom[19726] = 16'hffff;
  rom[19727] = 16'hdeda;
  rom[19728] = 16'h8bab;
  rom[19729] = 16'h7265;
  rom[19730] = 16'hb42a;
  rom[19731] = 16'he56d;
  rom[19732] = 16'hed6c;
  rom[19733] = 16'hfd8c;
  rom[19734] = 16'hf549;
  rom[19735] = 16'hfd68;
  rom[19736] = 16'hfd07;
  rom[19737] = 16'hfd27;
  rom[19738] = 16'hf508;
  rom[19739] = 16'hfd49;
  rom[19740] = 16'hf549;
  rom[19741] = 16'hed29;
  rom[19742] = 16'hf548;
  rom[19743] = 16'hecc6;
  rom[19744] = 16'hfd28;
  rom[19745] = 16'hfce8;
  rom[19746] = 16'hf54b;
  rom[19747] = 16'hdccb;
  rom[19748] = 16'h8b27;
  rom[19749] = 16'hc531;
  rom[19750] = 16'hfffe;
  rom[19751] = 16'hffff;
  rom[19752] = 16'hffff;
  rom[19753] = 16'hffff;
  rom[19754] = 16'hffff;
  rom[19755] = 16'hffff;
  rom[19756] = 16'hffff;
  rom[19757] = 16'hffff;
  rom[19758] = 16'hffff;
  rom[19759] = 16'hffff;
  rom[19760] = 16'hffff;
  rom[19761] = 16'hffff;
  rom[19762] = 16'hffff;
  rom[19763] = 16'hffff;
  rom[19764] = 16'hffff;
  rom[19765] = 16'hffff;
  rom[19766] = 16'hffff;
  rom[19767] = 16'hffff;
  rom[19768] = 16'hffff;
  rom[19769] = 16'hffff;
  rom[19770] = 16'hffff;
  rom[19771] = 16'hffff;
  rom[19772] = 16'hffff;
  rom[19773] = 16'hffff;
  rom[19774] = 16'hffff;
  rom[19775] = 16'hffff;
  rom[19776] = 16'hffff;
  rom[19777] = 16'hffff;
  rom[19778] = 16'hffff;
  rom[19779] = 16'hffff;
  rom[19780] = 16'hffff;
  rom[19781] = 16'hffff;
  rom[19782] = 16'hffff;
  rom[19783] = 16'hffff;
  rom[19784] = 16'hffff;
  rom[19785] = 16'hffff;
  rom[19786] = 16'hffff;
  rom[19787] = 16'hffff;
  rom[19788] = 16'hffff;
  rom[19789] = 16'hffff;
  rom[19790] = 16'hffff;
  rom[19791] = 16'hffff;
  rom[19792] = 16'hffff;
  rom[19793] = 16'hffff;
  rom[19794] = 16'hffff;
  rom[19795] = 16'hffff;
  rom[19796] = 16'hffff;
  rom[19797] = 16'hffff;
  rom[19798] = 16'hffff;
  rom[19799] = 16'hffff;
  rom[19800] = 16'hffff;
  rom[19801] = 16'hffff;
  rom[19802] = 16'hffff;
  rom[19803] = 16'hffff;
  rom[19804] = 16'hffff;
  rom[19805] = 16'hffff;
  rom[19806] = 16'hffff;
  rom[19807] = 16'hffff;
  rom[19808] = 16'hffff;
  rom[19809] = 16'hffff;
  rom[19810] = 16'hffff;
  rom[19811] = 16'hffff;
  rom[19812] = 16'hffff;
  rom[19813] = 16'hffff;
  rom[19814] = 16'hffff;
  rom[19815] = 16'hffff;
  rom[19816] = 16'hffff;
  rom[19817] = 16'hffff;
  rom[19818] = 16'hffff;
  rom[19819] = 16'hffff;
  rom[19820] = 16'hffff;
  rom[19821] = 16'hffff;
  rom[19822] = 16'hffff;
  rom[19823] = 16'hffff;
  rom[19824] = 16'hffff;
  rom[19825] = 16'hffff;
  rom[19826] = 16'hffff;
  rom[19827] = 16'hffff;
  rom[19828] = 16'he6d9;
  rom[19829] = 16'h6b26;
  rom[19830] = 16'h83c6;
  rom[19831] = 16'hcdec;
  rom[19832] = 16'heeae;
  rom[19833] = 16'hff2d;
  rom[19834] = 16'hf709;
  rom[19835] = 16'hf708;
  rom[19836] = 16'hff29;
  rom[19837] = 16'hf729;
  rom[19838] = 16'hff4a;
  rom[19839] = 16'hff28;
  rom[19840] = 16'hff29;
  rom[19841] = 16'hff28;
  rom[19842] = 16'hff29;
  rom[19843] = 16'hff28;
  rom[19844] = 16'hff29;
  rom[19845] = 16'hf728;
  rom[19846] = 16'hff49;
  rom[19847] = 16'hff49;
  rom[19848] = 16'hf72a;
  rom[19849] = 16'hff4a;
  rom[19850] = 16'hff4b;
  rom[19851] = 16'hcd88;
  rom[19852] = 16'h69e1;
  rom[19853] = 16'hc469;
  rom[19854] = 16'hed4b;
  rom[19855] = 16'hf529;
  rom[19856] = 16'hfd29;
  rom[19857] = 16'hfd27;
  rom[19858] = 16'hfd48;
  rom[19859] = 16'hfd27;
  rom[19860] = 16'hfd49;
  rom[19861] = 16'hfd29;
  rom[19862] = 16'hfd4a;
  rom[19863] = 16'hed4b;
  rom[19864] = 16'hedae;
  rom[19865] = 16'hac6b;
  rom[19866] = 16'h6aa7;
  rom[19867] = 16'hfffe;
  rom[19868] = 16'hffff;
  rom[19869] = 16'hffff;
  rom[19870] = 16'hffff;
  rom[19871] = 16'hffff;
  rom[19872] = 16'hffff;
  rom[19873] = 16'hffff;
  rom[19874] = 16'hffff;
  rom[19875] = 16'hffff;
  rom[19876] = 16'hffff;
  rom[19877] = 16'hffff;
  rom[19878] = 16'hffff;
  rom[19879] = 16'hffff;
  rom[19880] = 16'hffff;
  rom[19881] = 16'hffff;
  rom[19882] = 16'hffff;
  rom[19883] = 16'hffff;
  rom[19884] = 16'hffff;
  rom[19885] = 16'hffff;
  rom[19886] = 16'hffff;
  rom[19887] = 16'hffff;
  rom[19888] = 16'hffff;
  rom[19889] = 16'hffff;
  rom[19890] = 16'hffff;
  rom[19891] = 16'hffff;
  rom[19892] = 16'hffff;
  rom[19893] = 16'hffff;
  rom[19894] = 16'hc618;
  rom[19895] = 16'h6b6d;
  rom[19896] = 16'h41e8;
  rom[19897] = 16'h3986;
  rom[19898] = 16'h62ec;
  rom[19899] = 16'ha514;
  rom[19900] = 16'hffdf;
  rom[19901] = 16'hffdf;
  rom[19902] = 16'hffff;
  rom[19903] = 16'hffff;
  rom[19904] = 16'hffff;
  rom[19905] = 16'hffff;
  rom[19906] = 16'hffff;
  rom[19907] = 16'hffff;
  rom[19908] = 16'hffff;
  rom[19909] = 16'hffff;
  rom[19910] = 16'hffff;
  rom[19911] = 16'hffff;
  rom[19912] = 16'hffff;
  rom[19913] = 16'hffff;
  rom[19914] = 16'hffff;
  rom[19915] = 16'hffff;
  rom[19916] = 16'hffff;
  rom[19917] = 16'hffff;
  rom[19918] = 16'hffff;
  rom[19919] = 16'hffff;
  rom[19920] = 16'hffff;
  rom[19921] = 16'hffff;
  rom[19922] = 16'hffff;
  rom[19923] = 16'hffff;
  rom[19924] = 16'hffff;
  rom[19925] = 16'hffff;
  rom[19926] = 16'hffff;
  rom[19927] = 16'had32;
  rom[19928] = 16'h8328;
  rom[19929] = 16'hdd4e;
  rom[19930] = 16'hed4b;
  rom[19931] = 16'hf54a;
  rom[19932] = 16'hf54a;
  rom[19933] = 16'hf529;
  rom[19934] = 16'hfd6a;
  rom[19935] = 16'hfd28;
  rom[19936] = 16'hfd28;
  rom[19937] = 16'hfd28;
  rom[19938] = 16'hfd28;
  rom[19939] = 16'hf528;
  rom[19940] = 16'hf549;
  rom[19941] = 16'hfd48;
  rom[19942] = 16'hfd28;
  rom[19943] = 16'hfd48;
  rom[19944] = 16'hfd29;
  rom[19945] = 16'hed2a;
  rom[19946] = 16'hdd0c;
  rom[19947] = 16'ha3a9;
  rom[19948] = 16'h93ab;
  rom[19949] = 16'hf75b;
  rom[19950] = 16'hffff;
  rom[19951] = 16'hffff;
  rom[19952] = 16'hffff;
  rom[19953] = 16'hffff;
  rom[19954] = 16'hffff;
  rom[19955] = 16'hffff;
  rom[19956] = 16'hffff;
  rom[19957] = 16'hffff;
  rom[19958] = 16'hffff;
  rom[19959] = 16'hffff;
  rom[19960] = 16'hffff;
  rom[19961] = 16'hffff;
  rom[19962] = 16'hffff;
  rom[19963] = 16'hffff;
  rom[19964] = 16'hffff;
  rom[19965] = 16'hffff;
  rom[19966] = 16'hffff;
  rom[19967] = 16'hffff;
  rom[19968] = 16'hffff;
  rom[19969] = 16'hffff;
  rom[19970] = 16'hffff;
  rom[19971] = 16'hffff;
  rom[19972] = 16'hffff;
  rom[19973] = 16'hffff;
  rom[19974] = 16'hffff;
  rom[19975] = 16'hffff;
  rom[19976] = 16'hffff;
  rom[19977] = 16'hffff;
  rom[19978] = 16'hffff;
  rom[19979] = 16'hffff;
  rom[19980] = 16'hffff;
  rom[19981] = 16'hffff;
  rom[19982] = 16'hffff;
  rom[19983] = 16'hffff;
  rom[19984] = 16'hffff;
  rom[19985] = 16'hffff;
  rom[19986] = 16'hffff;
  rom[19987] = 16'hffff;
  rom[19988] = 16'hffff;
  rom[19989] = 16'hffff;
  rom[19990] = 16'hffff;
  rom[19991] = 16'hffff;
  rom[19992] = 16'hffff;
  rom[19993] = 16'hffff;
  rom[19994] = 16'hffff;
  rom[19995] = 16'hffff;
  rom[19996] = 16'hffff;
  rom[19997] = 16'hffff;
  rom[19998] = 16'hffff;
  rom[19999] = 16'hffff;
  rom[20000] = 16'hffff;
  rom[20001] = 16'hffff;
  rom[20002] = 16'hffff;
  rom[20003] = 16'hffff;
  rom[20004] = 16'hffff;
  rom[20005] = 16'hffff;
  rom[20006] = 16'hffff;
  rom[20007] = 16'hffff;
  rom[20008] = 16'hffff;
  rom[20009] = 16'hffff;
  rom[20010] = 16'hffff;
  rom[20011] = 16'hffff;
  rom[20012] = 16'hffff;
  rom[20013] = 16'hffff;
  rom[20014] = 16'hffff;
  rom[20015] = 16'hffff;
  rom[20016] = 16'hffff;
  rom[20017] = 16'hffff;
  rom[20018] = 16'hffff;
  rom[20019] = 16'hffff;
  rom[20020] = 16'hffff;
  rom[20021] = 16'hffff;
  rom[20022] = 16'hffff;
  rom[20023] = 16'hffff;
  rom[20024] = 16'hffde;
  rom[20025] = 16'hffff;
  rom[20026] = 16'hffff;
  rom[20027] = 16'hffdf;
  rom[20028] = 16'hfffe;
  rom[20029] = 16'hded8;
  rom[20030] = 16'h7348;
  rom[20031] = 16'h5241;
  rom[20032] = 16'h9447;
  rom[20033] = 16'heece;
  rom[20034] = 16'hff6b;
  rom[20035] = 16'hff29;
  rom[20036] = 16'hf709;
  rom[20037] = 16'hff29;
  rom[20038] = 16'hf6e8;
  rom[20039] = 16'hff29;
  rom[20040] = 16'hf708;
  rom[20041] = 16'hff28;
  rom[20042] = 16'hff08;
  rom[20043] = 16'hff28;
  rom[20044] = 16'hf708;
  rom[20045] = 16'hf729;
  rom[20046] = 16'hf728;
  rom[20047] = 16'hff49;
  rom[20048] = 16'hf709;
  rom[20049] = 16'hf70a;
  rom[20050] = 16'hf6e9;
  rom[20051] = 16'hfeea;
  rom[20052] = 16'h7ac1;
  rom[20053] = 16'h7a63;
  rom[20054] = 16'he50a;
  rom[20055] = 16'hece9;
  rom[20056] = 16'hf549;
  rom[20057] = 16'hfd48;
  rom[20058] = 16'hf506;
  rom[20059] = 16'hf527;
  rom[20060] = 16'hf548;
  rom[20061] = 16'hfd28;
  rom[20062] = 16'hfd28;
  rom[20063] = 16'hfd49;
  rom[20064] = 16'he509;
  rom[20065] = 16'hc4ec;
  rom[20066] = 16'h838a;
  rom[20067] = 16'hffff;
  rom[20068] = 16'hf7ff;
  rom[20069] = 16'hffff;
  rom[20070] = 16'hffff;
  rom[20071] = 16'hffff;
  rom[20072] = 16'hffff;
  rom[20073] = 16'hffff;
  rom[20074] = 16'hffff;
  rom[20075] = 16'hffff;
  rom[20076] = 16'hffff;
  rom[20077] = 16'hffff;
  rom[20078] = 16'hffff;
  rom[20079] = 16'hffff;
  rom[20080] = 16'hffff;
  rom[20081] = 16'hffff;
  rom[20082] = 16'hffdf;
  rom[20083] = 16'hffff;
  rom[20084] = 16'hffff;
  rom[20085] = 16'hffff;
  rom[20086] = 16'hffff;
  rom[20087] = 16'hffff;
  rom[20088] = 16'hffff;
  rom[20089] = 16'hffff;
  rom[20090] = 16'hffff;
  rom[20091] = 16'hffff;
  rom[20092] = 16'hffff;
  rom[20093] = 16'hb596;
  rom[20094] = 16'h39c6;
  rom[20095] = 16'h41c7;
  rom[20096] = 16'h8c30;
  rom[20097] = 16'h9492;
  rom[20098] = 16'h528a;
  rom[20099] = 16'h41c7;
  rom[20100] = 16'h9451;
  rom[20101] = 16'hffbf;
  rom[20102] = 16'hffff;
  rom[20103] = 16'hffff;
  rom[20104] = 16'hffff;
  rom[20105] = 16'hffff;
  rom[20106] = 16'hffff;
  rom[20107] = 16'hffff;
  rom[20108] = 16'hffff;
  rom[20109] = 16'hffff;
  rom[20110] = 16'hffff;
  rom[20111] = 16'hffff;
  rom[20112] = 16'hffff;
  rom[20113] = 16'hffff;
  rom[20114] = 16'hffff;
  rom[20115] = 16'hffff;
  rom[20116] = 16'hffff;
  rom[20117] = 16'hffff;
  rom[20118] = 16'hffff;
  rom[20119] = 16'hffff;
  rom[20120] = 16'hffff;
  rom[20121] = 16'hffff;
  rom[20122] = 16'hffff;
  rom[20123] = 16'hffff;
  rom[20124] = 16'hffff;
  rom[20125] = 16'hffff;
  rom[20126] = 16'hf7be;
  rom[20127] = 16'hc5f5;
  rom[20128] = 16'h93a8;
  rom[20129] = 16'hdd0a;
  rom[20130] = 16'hf548;
  rom[20131] = 16'hfd88;
  rom[20132] = 16'hfd27;
  rom[20133] = 16'hfd28;
  rom[20134] = 16'hf4e7;
  rom[20135] = 16'hfd28;
  rom[20136] = 16'hf508;
  rom[20137] = 16'hfd28;
  rom[20138] = 16'hfd28;
  rom[20139] = 16'hfd48;
  rom[20140] = 16'hf527;
  rom[20141] = 16'hf507;
  rom[20142] = 16'hfd48;
  rom[20143] = 16'hf4e7;
  rom[20144] = 16'hece8;
  rom[20145] = 16'hf5ad;
  rom[20146] = 16'hb46b;
  rom[20147] = 16'h6a87;
  rom[20148] = 16'hd677;
  rom[20149] = 16'hffff;
  rom[20150] = 16'hffff;
  rom[20151] = 16'hffff;
  rom[20152] = 16'hffff;
  rom[20153] = 16'hffff;
  rom[20154] = 16'hffff;
  rom[20155] = 16'hffff;
  rom[20156] = 16'hffff;
  rom[20157] = 16'hffff;
  rom[20158] = 16'hffff;
  rom[20159] = 16'hffff;
  rom[20160] = 16'hffff;
  rom[20161] = 16'hffff;
  rom[20162] = 16'hffff;
  rom[20163] = 16'hffff;
  rom[20164] = 16'hffff;
  rom[20165] = 16'hffff;
  rom[20166] = 16'hffff;
  rom[20167] = 16'hffff;
  rom[20168] = 16'hffff;
  rom[20169] = 16'hffff;
  rom[20170] = 16'hffff;
  rom[20171] = 16'hffff;
  rom[20172] = 16'hffff;
  rom[20173] = 16'hffff;
  rom[20174] = 16'hffff;
  rom[20175] = 16'hffff;
  rom[20176] = 16'hffff;
  rom[20177] = 16'hffff;
  rom[20178] = 16'hffff;
  rom[20179] = 16'hffff;
  rom[20180] = 16'hffff;
  rom[20181] = 16'hffff;
  rom[20182] = 16'hffff;
  rom[20183] = 16'hffff;
  rom[20184] = 16'hffff;
  rom[20185] = 16'hffff;
  rom[20186] = 16'hffff;
  rom[20187] = 16'hffff;
  rom[20188] = 16'hffff;
  rom[20189] = 16'hffff;
  rom[20190] = 16'hffff;
  rom[20191] = 16'hffff;
  rom[20192] = 16'hffff;
  rom[20193] = 16'hffff;
  rom[20194] = 16'hffff;
  rom[20195] = 16'hffff;
  rom[20196] = 16'hffff;
  rom[20197] = 16'hffff;
  rom[20198] = 16'hffff;
  rom[20199] = 16'hffff;
  rom[20200] = 16'hffff;
  rom[20201] = 16'hffff;
  rom[20202] = 16'hffff;
  rom[20203] = 16'hffff;
  rom[20204] = 16'hffff;
  rom[20205] = 16'hffff;
  rom[20206] = 16'hffff;
  rom[20207] = 16'hffff;
  rom[20208] = 16'hffff;
  rom[20209] = 16'hffff;
  rom[20210] = 16'hffff;
  rom[20211] = 16'hffff;
  rom[20212] = 16'hffff;
  rom[20213] = 16'hffff;
  rom[20214] = 16'hffff;
  rom[20215] = 16'hffff;
  rom[20216] = 16'hffff;
  rom[20217] = 16'hffff;
  rom[20218] = 16'hffff;
  rom[20219] = 16'hffff;
  rom[20220] = 16'hffff;
  rom[20221] = 16'hffff;
  rom[20222] = 16'hffff;
  rom[20223] = 16'hffff;
  rom[20224] = 16'hffff;
  rom[20225] = 16'hffff;
  rom[20226] = 16'hffff;
  rom[20227] = 16'hffff;
  rom[20228] = 16'hffff;
  rom[20229] = 16'hffff;
  rom[20230] = 16'hf77c;
  rom[20231] = 16'hb571;
  rom[20232] = 16'h7346;
  rom[20233] = 16'hbdac;
  rom[20234] = 16'hf72c;
  rom[20235] = 16'hf72a;
  rom[20236] = 16'hf729;
  rom[20237] = 16'hf728;
  rom[20238] = 16'hff49;
  rom[20239] = 16'hff29;
  rom[20240] = 16'hff2a;
  rom[20241] = 16'hf729;
  rom[20242] = 16'hff49;
  rom[20243] = 16'hff28;
  rom[20244] = 16'hff2a;
  rom[20245] = 16'hf72a;
  rom[20246] = 16'hff2a;
  rom[20247] = 16'hff2a;
  rom[20248] = 16'hff0a;
  rom[20249] = 16'hf729;
  rom[20250] = 16'hff29;
  rom[20251] = 16'hf70a;
  rom[20252] = 16'he5eb;
  rom[20253] = 16'h6a00;
  rom[20254] = 16'hcc68;
  rom[20255] = 16'hed0a;
  rom[20256] = 16'hf56a;
  rom[20257] = 16'hf507;
  rom[20258] = 16'hfd47;
  rom[20259] = 16'hfd47;
  rom[20260] = 16'hfd27;
  rom[20261] = 16'hfd27;
  rom[20262] = 16'hfd28;
  rom[20263] = 16'hfd28;
  rom[20264] = 16'hed4a;
  rom[20265] = 16'hc4cb;
  rom[20266] = 16'ha44d;
  rom[20267] = 16'hfffe;
  rom[20268] = 16'hffff;
  rom[20269] = 16'hffff;
  rom[20270] = 16'hffff;
  rom[20271] = 16'hffff;
  rom[20272] = 16'hffff;
  rom[20273] = 16'hffff;
  rom[20274] = 16'hffff;
  rom[20275] = 16'hffff;
  rom[20276] = 16'hffff;
  rom[20277] = 16'hffff;
  rom[20278] = 16'hffff;
  rom[20279] = 16'hffff;
  rom[20280] = 16'hffff;
  rom[20281] = 16'hffff;
  rom[20282] = 16'hffff;
  rom[20283] = 16'hffff;
  rom[20284] = 16'hffff;
  rom[20285] = 16'hffff;
  rom[20286] = 16'hffff;
  rom[20287] = 16'hffff;
  rom[20288] = 16'hffff;
  rom[20289] = 16'hffff;
  rom[20290] = 16'hffff;
  rom[20291] = 16'hffff;
  rom[20292] = 16'hef5d;
  rom[20293] = 16'h5289;
  rom[20294] = 16'h62cb;
  rom[20295] = 16'hde9a;
  rom[20296] = 16'hffff;
  rom[20297] = 16'hffbe;
  rom[20298] = 16'hff5e;
  rom[20299] = 16'h7b8e;
  rom[20300] = 16'h41c7;
  rom[20301] = 16'hc5f8;
  rom[20302] = 16'hffff;
  rom[20303] = 16'hffff;
  rom[20304] = 16'hffff;
  rom[20305] = 16'hffff;
  rom[20306] = 16'hffff;
  rom[20307] = 16'hffff;
  rom[20308] = 16'hffff;
  rom[20309] = 16'hffff;
  rom[20310] = 16'hffff;
  rom[20311] = 16'hffff;
  rom[20312] = 16'hffff;
  rom[20313] = 16'hffff;
  rom[20314] = 16'hffff;
  rom[20315] = 16'hffff;
  rom[20316] = 16'hffff;
  rom[20317] = 16'hffff;
  rom[20318] = 16'hffff;
  rom[20319] = 16'hffff;
  rom[20320] = 16'hffff;
  rom[20321] = 16'hffff;
  rom[20322] = 16'hffff;
  rom[20323] = 16'hffff;
  rom[20324] = 16'hffff;
  rom[20325] = 16'hffff;
  rom[20326] = 16'hffff;
  rom[20327] = 16'hce14;
  rom[20328] = 16'h9388;
  rom[20329] = 16'he54b;
  rom[20330] = 16'hfd49;
  rom[20331] = 16'hf4e5;
  rom[20332] = 16'hfd67;
  rom[20333] = 16'hfd07;
  rom[20334] = 16'hfd4a;
  rom[20335] = 16'hfd09;
  rom[20336] = 16'hfd49;
  rom[20337] = 16'hf527;
  rom[20338] = 16'hfd28;
  rom[20339] = 16'hf528;
  rom[20340] = 16'hfd28;
  rom[20341] = 16'hfd27;
  rom[20342] = 16'hfd28;
  rom[20343] = 16'hf4e7;
  rom[20344] = 16'hf56b;
  rom[20345] = 16'hd4ec;
  rom[20346] = 16'h7ae8;
  rom[20347] = 16'hbdb4;
  rom[20348] = 16'hffff;
  rom[20349] = 16'hffdf;
  rom[20350] = 16'hffff;
  rom[20351] = 16'hffff;
  rom[20352] = 16'hffff;
  rom[20353] = 16'hffff;
  rom[20354] = 16'hffff;
  rom[20355] = 16'hffff;
  rom[20356] = 16'hffff;
  rom[20357] = 16'hffff;
  rom[20358] = 16'hffff;
  rom[20359] = 16'hffff;
  rom[20360] = 16'hffff;
  rom[20361] = 16'hffff;
  rom[20362] = 16'hffff;
  rom[20363] = 16'hffff;
  rom[20364] = 16'hffff;
  rom[20365] = 16'hffff;
  rom[20366] = 16'hffff;
  rom[20367] = 16'hffff;
  rom[20368] = 16'hffff;
  rom[20369] = 16'hffff;
  rom[20370] = 16'hffff;
  rom[20371] = 16'hffff;
  rom[20372] = 16'hffff;
  rom[20373] = 16'hffff;
  rom[20374] = 16'hffff;
  rom[20375] = 16'hffff;
  rom[20376] = 16'hffff;
  rom[20377] = 16'hffff;
  rom[20378] = 16'hffff;
  rom[20379] = 16'hffff;
  rom[20380] = 16'hffff;
  rom[20381] = 16'hffff;
  rom[20382] = 16'hffff;
  rom[20383] = 16'hffff;
  rom[20384] = 16'hffff;
  rom[20385] = 16'hffff;
  rom[20386] = 16'hffff;
  rom[20387] = 16'hffff;
  rom[20388] = 16'hffff;
  rom[20389] = 16'hffff;
  rom[20390] = 16'hffff;
  rom[20391] = 16'hffff;
  rom[20392] = 16'hffff;
  rom[20393] = 16'hffff;
  rom[20394] = 16'hffff;
  rom[20395] = 16'hffff;
  rom[20396] = 16'hffff;
  rom[20397] = 16'hffff;
  rom[20398] = 16'hffff;
  rom[20399] = 16'hffff;
  rom[20400] = 16'hffff;
  rom[20401] = 16'hffff;
  rom[20402] = 16'hffff;
  rom[20403] = 16'hffff;
  rom[20404] = 16'hffff;
  rom[20405] = 16'hffff;
  rom[20406] = 16'hffff;
  rom[20407] = 16'hffff;
  rom[20408] = 16'hffff;
  rom[20409] = 16'hffff;
  rom[20410] = 16'hffff;
  rom[20411] = 16'hffff;
  rom[20412] = 16'hffff;
  rom[20413] = 16'hffff;
  rom[20414] = 16'hffff;
  rom[20415] = 16'hffff;
  rom[20416] = 16'hffff;
  rom[20417] = 16'hffff;
  rom[20418] = 16'hffff;
  rom[20419] = 16'hffff;
  rom[20420] = 16'hffff;
  rom[20421] = 16'hffff;
  rom[20422] = 16'hffff;
  rom[20423] = 16'hffff;
  rom[20424] = 16'hffbf;
  rom[20425] = 16'hffff;
  rom[20426] = 16'hffdf;
  rom[20427] = 16'hffff;
  rom[20428] = 16'hffff;
  rom[20429] = 16'hffff;
  rom[20430] = 16'hffdf;
  rom[20431] = 16'hffbd;
  rom[20432] = 16'h944c;
  rom[20433] = 16'h7365;
  rom[20434] = 16'he6cd;
  rom[20435] = 16'hff6c;
  rom[20436] = 16'hf709;
  rom[20437] = 16'hff48;
  rom[20438] = 16'hf708;
  rom[20439] = 16'hff2a;
  rom[20440] = 16'hf72a;
  rom[20441] = 16'hf729;
  rom[20442] = 16'hf728;
  rom[20443] = 16'hff28;
  rom[20444] = 16'hfee9;
  rom[20445] = 16'hff29;
  rom[20446] = 16'hf709;
  rom[20447] = 16'hff0a;
  rom[20448] = 16'hff09;
  rom[20449] = 16'hff29;
  rom[20450] = 16'hf729;
  rom[20451] = 16'hf72a;
  rom[20452] = 16'hff0d;
  rom[20453] = 16'ha405;
  rom[20454] = 16'h8ac2;
  rom[20455] = 16'he50a;
  rom[20456] = 16'hed09;
  rom[20457] = 16'hfd68;
  rom[20458] = 16'hfd27;
  rom[20459] = 16'hfd27;
  rom[20460] = 16'hfd07;
  rom[20461] = 16'hfd28;
  rom[20462] = 16'hfd08;
  rom[20463] = 16'hfd4a;
  rom[20464] = 16'hed4b;
  rom[20465] = 16'hc48b;
  rom[20466] = 16'hacae;
  rom[20467] = 16'hffdd;
  rom[20468] = 16'hffff;
  rom[20469] = 16'hffff;
  rom[20470] = 16'hffff;
  rom[20471] = 16'hffff;
  rom[20472] = 16'hffff;
  rom[20473] = 16'hffff;
  rom[20474] = 16'hffff;
  rom[20475] = 16'hffff;
  rom[20476] = 16'hffff;
  rom[20477] = 16'hffff;
  rom[20478] = 16'hffff;
  rom[20479] = 16'hffff;
  rom[20480] = 16'hffff;
  rom[20481] = 16'hffff;
  rom[20482] = 16'hffff;
  rom[20483] = 16'hffff;
  rom[20484] = 16'hffff;
  rom[20485] = 16'hffff;
  rom[20486] = 16'hffff;
  rom[20487] = 16'hffff;
  rom[20488] = 16'hffff;
  rom[20489] = 16'hffff;
  rom[20490] = 16'hffff;
  rom[20491] = 16'hffff;
  rom[20492] = 16'ha534;
  rom[20493] = 16'h2103;
  rom[20494] = 16'hbd96;
  rom[20495] = 16'hffff;
  rom[20496] = 16'hffff;
  rom[20497] = 16'hffbf;
  rom[20498] = 16'hffdf;
  rom[20499] = 16'he6dc;
  rom[20500] = 16'h4a48;
  rom[20501] = 16'h83cf;
  rom[20502] = 16'hff7e;
  rom[20503] = 16'hffff;
  rom[20504] = 16'hffff;
  rom[20505] = 16'hffff;
  rom[20506] = 16'hffff;
  rom[20507] = 16'hffff;
  rom[20508] = 16'hffff;
  rom[20509] = 16'hffff;
  rom[20510] = 16'hffff;
  rom[20511] = 16'hffff;
  rom[20512] = 16'hffff;
  rom[20513] = 16'hffff;
  rom[20514] = 16'hffff;
  rom[20515] = 16'hffff;
  rom[20516] = 16'hffff;
  rom[20517] = 16'hffff;
  rom[20518] = 16'hffff;
  rom[20519] = 16'hffff;
  rom[20520] = 16'hffff;
  rom[20521] = 16'hffff;
  rom[20522] = 16'hffff;
  rom[20523] = 16'hffff;
  rom[20524] = 16'hffdf;
  rom[20525] = 16'hffff;
  rom[20526] = 16'hffff;
  rom[20527] = 16'hd676;
  rom[20528] = 16'h8b67;
  rom[20529] = 16'hdceb;
  rom[20530] = 16'hf549;
  rom[20531] = 16'hfd27;
  rom[20532] = 16'hf526;
  rom[20533] = 16'hfd48;
  rom[20534] = 16'hf508;
  rom[20535] = 16'hfd29;
  rom[20536] = 16'hfce8;
  rom[20537] = 16'hfd48;
  rom[20538] = 16'hf507;
  rom[20539] = 16'hfd49;
  rom[20540] = 16'hfd29;
  rom[20541] = 16'hfd28;
  rom[20542] = 16'hf507;
  rom[20543] = 16'hece8;
  rom[20544] = 16'hdd0b;
  rom[20545] = 16'h8aa5;
  rom[20546] = 16'h9c4e;
  rom[20547] = 16'hf7be;
  rom[20548] = 16'hffff;
  rom[20549] = 16'hffff;
  rom[20550] = 16'hffff;
  rom[20551] = 16'hffff;
  rom[20552] = 16'hffff;
  rom[20553] = 16'hffff;
  rom[20554] = 16'hffff;
  rom[20555] = 16'hffff;
  rom[20556] = 16'hffff;
  rom[20557] = 16'hffff;
  rom[20558] = 16'hffff;
  rom[20559] = 16'hffff;
  rom[20560] = 16'hffff;
  rom[20561] = 16'hffff;
  rom[20562] = 16'hffff;
  rom[20563] = 16'hffff;
  rom[20564] = 16'hffff;
  rom[20565] = 16'hffff;
  rom[20566] = 16'hffff;
  rom[20567] = 16'hffff;
  rom[20568] = 16'hffff;
  rom[20569] = 16'hffff;
  rom[20570] = 16'hffff;
  rom[20571] = 16'hffff;
  rom[20572] = 16'hffff;
  rom[20573] = 16'hffff;
  rom[20574] = 16'hffff;
  rom[20575] = 16'hffff;
  rom[20576] = 16'hffff;
  rom[20577] = 16'hffff;
  rom[20578] = 16'hffff;
  rom[20579] = 16'hffff;
  rom[20580] = 16'hffff;
  rom[20581] = 16'hffff;
  rom[20582] = 16'hffff;
  rom[20583] = 16'hffff;
  rom[20584] = 16'hffff;
  rom[20585] = 16'hffff;
  rom[20586] = 16'hffff;
  rom[20587] = 16'hffff;
  rom[20588] = 16'hffff;
  rom[20589] = 16'hffff;
  rom[20590] = 16'hffff;
  rom[20591] = 16'hffff;
  rom[20592] = 16'hffff;
  rom[20593] = 16'hffff;
  rom[20594] = 16'hffff;
  rom[20595] = 16'hffff;
  rom[20596] = 16'hffff;
  rom[20597] = 16'hffff;
  rom[20598] = 16'hffff;
  rom[20599] = 16'hffff;
  rom[20600] = 16'hffff;
  rom[20601] = 16'hffff;
  rom[20602] = 16'hffff;
  rom[20603] = 16'hffff;
  rom[20604] = 16'hffff;
  rom[20605] = 16'hffff;
  rom[20606] = 16'hffff;
  rom[20607] = 16'hffff;
  rom[20608] = 16'hffff;
  rom[20609] = 16'hffff;
  rom[20610] = 16'hffff;
  rom[20611] = 16'hffff;
  rom[20612] = 16'hffff;
  rom[20613] = 16'hffff;
  rom[20614] = 16'hffff;
  rom[20615] = 16'hffff;
  rom[20616] = 16'hffff;
  rom[20617] = 16'hffff;
  rom[20618] = 16'hffff;
  rom[20619] = 16'hffff;
  rom[20620] = 16'hffff;
  rom[20621] = 16'hffff;
  rom[20622] = 16'hffff;
  rom[20623] = 16'hffff;
  rom[20624] = 16'hffff;
  rom[20625] = 16'hffff;
  rom[20626] = 16'hffff;
  rom[20627] = 16'hffff;
  rom[20628] = 16'hffff;
  rom[20629] = 16'hffff;
  rom[20630] = 16'hffff;
  rom[20631] = 16'hffde;
  rom[20632] = 16'heef9;
  rom[20633] = 16'h6b05;
  rom[20634] = 16'h9c87;
  rom[20635] = 16'he6cb;
  rom[20636] = 16'hf70a;
  rom[20637] = 16'hff29;
  rom[20638] = 16'hff2a;
  rom[20639] = 16'hf70b;
  rom[20640] = 16'hf74b;
  rom[20641] = 16'hf749;
  rom[20642] = 16'hf748;
  rom[20643] = 16'hff48;
  rom[20644] = 16'hff49;
  rom[20645] = 16'hff29;
  rom[20646] = 16'hff29;
  rom[20647] = 16'hff09;
  rom[20648] = 16'hff2a;
  rom[20649] = 16'hff28;
  rom[20650] = 16'hf74a;
  rom[20651] = 16'hf70a;
  rom[20652] = 16'hf70c;
  rom[20653] = 16'hddca;
  rom[20654] = 16'h7a42;
  rom[20655] = 16'hc408;
  rom[20656] = 16'hf54c;
  rom[20657] = 16'hf529;
  rom[20658] = 16'hfd28;
  rom[20659] = 16'hfce7;
  rom[20660] = 16'hfd28;
  rom[20661] = 16'hfd29;
  rom[20662] = 16'hfd29;
  rom[20663] = 16'hf528;
  rom[20664] = 16'hf5ac;
  rom[20665] = 16'hbc8a;
  rom[20666] = 16'hb4ad;
  rom[20667] = 16'hfffd;
  rom[20668] = 16'hffff;
  rom[20669] = 16'hffff;
  rom[20670] = 16'hffff;
  rom[20671] = 16'hffff;
  rom[20672] = 16'hffff;
  rom[20673] = 16'hffff;
  rom[20674] = 16'hffff;
  rom[20675] = 16'hffff;
  rom[20676] = 16'hffff;
  rom[20677] = 16'hffff;
  rom[20678] = 16'hffff;
  rom[20679] = 16'hffff;
  rom[20680] = 16'hffff;
  rom[20681] = 16'hffff;
  rom[20682] = 16'hffff;
  rom[20683] = 16'hffff;
  rom[20684] = 16'hffff;
  rom[20685] = 16'hffff;
  rom[20686] = 16'hffff;
  rom[20687] = 16'hffff;
  rom[20688] = 16'hffff;
  rom[20689] = 16'hffff;
  rom[20690] = 16'hffff;
  rom[20691] = 16'hffff;
  rom[20692] = 16'hce39;
  rom[20693] = 16'h9472;
  rom[20694] = 16'hf79e;
  rom[20695] = 16'hf7bf;
  rom[20696] = 16'hffff;
  rom[20697] = 16'hffff;
  rom[20698] = 16'hffff;
  rom[20699] = 16'hffff;
  rom[20700] = 16'hbdb7;
  rom[20701] = 16'hb5b6;
  rom[20702] = 16'hffff;
  rom[20703] = 16'hffff;
  rom[20704] = 16'hffff;
  rom[20705] = 16'hffff;
  rom[20706] = 16'hffff;
  rom[20707] = 16'hffff;
  rom[20708] = 16'hffff;
  rom[20709] = 16'hffff;
  rom[20710] = 16'hffff;
  rom[20711] = 16'hffff;
  rom[20712] = 16'hffff;
  rom[20713] = 16'hffff;
  rom[20714] = 16'hffff;
  rom[20715] = 16'hffff;
  rom[20716] = 16'hffff;
  rom[20717] = 16'hffff;
  rom[20718] = 16'hffff;
  rom[20719] = 16'hffff;
  rom[20720] = 16'hffff;
  rom[20721] = 16'hffff;
  rom[20722] = 16'hffff;
  rom[20723] = 16'hffff;
  rom[20724] = 16'hffff;
  rom[20725] = 16'hffff;
  rom[20726] = 16'hffff;
  rom[20727] = 16'hd656;
  rom[20728] = 16'h9368;
  rom[20729] = 16'hed6d;
  rom[20730] = 16'hfd49;
  rom[20731] = 16'hfd27;
  rom[20732] = 16'hfd67;
  rom[20733] = 16'hfd27;
  rom[20734] = 16'hfd29;
  rom[20735] = 16'hfd29;
  rom[20736] = 16'hfd08;
  rom[20737] = 16'hf528;
  rom[20738] = 16'hfd6a;
  rom[20739] = 16'hed28;
  rom[20740] = 16'hf52a;
  rom[20741] = 16'hf509;
  rom[20742] = 16'hf52a;
  rom[20743] = 16'he54b;
  rom[20744] = 16'h9346;
  rom[20745] = 16'ha44d;
  rom[20746] = 16'hffbd;
  rom[20747] = 16'hffff;
  rom[20748] = 16'hffff;
  rom[20749] = 16'hffff;
  rom[20750] = 16'hffff;
  rom[20751] = 16'hffff;
  rom[20752] = 16'hffff;
  rom[20753] = 16'hffff;
  rom[20754] = 16'hffff;
  rom[20755] = 16'hffff;
  rom[20756] = 16'hffff;
  rom[20757] = 16'hffff;
  rom[20758] = 16'hffff;
  rom[20759] = 16'hffff;
  rom[20760] = 16'hffff;
  rom[20761] = 16'hffff;
  rom[20762] = 16'hffff;
  rom[20763] = 16'hffff;
  rom[20764] = 16'hffff;
  rom[20765] = 16'hffff;
  rom[20766] = 16'hffff;
  rom[20767] = 16'hffff;
  rom[20768] = 16'hffff;
  rom[20769] = 16'hffff;
  rom[20770] = 16'hffff;
  rom[20771] = 16'hffff;
  rom[20772] = 16'hffff;
  rom[20773] = 16'hffff;
  rom[20774] = 16'hffff;
  rom[20775] = 16'hffff;
  rom[20776] = 16'hffff;
  rom[20777] = 16'hffff;
  rom[20778] = 16'hffff;
  rom[20779] = 16'hffff;
  rom[20780] = 16'hffff;
  rom[20781] = 16'hffff;
  rom[20782] = 16'hffff;
  rom[20783] = 16'hffff;
  rom[20784] = 16'hffff;
  rom[20785] = 16'hffff;
  rom[20786] = 16'hffff;
  rom[20787] = 16'hffff;
  rom[20788] = 16'hffff;
  rom[20789] = 16'hffff;
  rom[20790] = 16'hffff;
  rom[20791] = 16'hffff;
  rom[20792] = 16'hffff;
  rom[20793] = 16'hffff;
  rom[20794] = 16'hffff;
  rom[20795] = 16'hffff;
  rom[20796] = 16'hffff;
  rom[20797] = 16'hffff;
  rom[20798] = 16'hffff;
  rom[20799] = 16'hffff;
  rom[20800] = 16'hffff;
  rom[20801] = 16'hffff;
  rom[20802] = 16'hffff;
  rom[20803] = 16'hffff;
  rom[20804] = 16'hffff;
  rom[20805] = 16'hffff;
  rom[20806] = 16'hffff;
  rom[20807] = 16'hffff;
  rom[20808] = 16'hffff;
  rom[20809] = 16'hffff;
  rom[20810] = 16'hffff;
  rom[20811] = 16'hffff;
  rom[20812] = 16'hffff;
  rom[20813] = 16'hffff;
  rom[20814] = 16'hffff;
  rom[20815] = 16'hffff;
  rom[20816] = 16'hffff;
  rom[20817] = 16'hffff;
  rom[20818] = 16'hffff;
  rom[20819] = 16'hffff;
  rom[20820] = 16'hffff;
  rom[20821] = 16'hffff;
  rom[20822] = 16'hffff;
  rom[20823] = 16'hffff;
  rom[20824] = 16'hffff;
  rom[20825] = 16'hffff;
  rom[20826] = 16'hffff;
  rom[20827] = 16'hffff;
  rom[20828] = 16'hffff;
  rom[20829] = 16'hffff;
  rom[20830] = 16'hffff;
  rom[20831] = 16'hffff;
  rom[20832] = 16'hfffd;
  rom[20833] = 16'hb551;
  rom[20834] = 16'h6b04;
  rom[20835] = 16'hc5cb;
  rom[20836] = 16'hef0c;
  rom[20837] = 16'hff2b;
  rom[20838] = 16'hf70b;
  rom[20839] = 16'hff0a;
  rom[20840] = 16'hf749;
  rom[20841] = 16'hef28;
  rom[20842] = 16'hf748;
  rom[20843] = 16'hf748;
  rom[20844] = 16'hf728;
  rom[20845] = 16'hff48;
  rom[20846] = 16'hff08;
  rom[20847] = 16'hff29;
  rom[20848] = 16'hf709;
  rom[20849] = 16'hff28;
  rom[20850] = 16'hf729;
  rom[20851] = 16'hff2a;
  rom[20852] = 16'hf70a;
  rom[20853] = 16'hf6ad;
  rom[20854] = 16'hac05;
  rom[20855] = 16'h7a21;
  rom[20856] = 16'hdcca;
  rom[20857] = 16'hed0a;
  rom[20858] = 16'hfd29;
  rom[20859] = 16'hfd29;
  rom[20860] = 16'hfd29;
  rom[20861] = 16'hfd29;
  rom[20862] = 16'hfd08;
  rom[20863] = 16'hfd49;
  rom[20864] = 16'he509;
  rom[20865] = 16'hccca;
  rom[20866] = 16'hac6b;
  rom[20867] = 16'hfffd;
  rom[20868] = 16'hffff;
  rom[20869] = 16'hffff;
  rom[20870] = 16'hffff;
  rom[20871] = 16'hffff;
  rom[20872] = 16'hffff;
  rom[20873] = 16'hffff;
  rom[20874] = 16'hffff;
  rom[20875] = 16'hffff;
  rom[20876] = 16'hffff;
  rom[20877] = 16'hffff;
  rom[20878] = 16'hffff;
  rom[20879] = 16'hffff;
  rom[20880] = 16'hffff;
  rom[20881] = 16'hffff;
  rom[20882] = 16'hffff;
  rom[20883] = 16'hffff;
  rom[20884] = 16'hffff;
  rom[20885] = 16'hffff;
  rom[20886] = 16'hffdf;
  rom[20887] = 16'hffff;
  rom[20888] = 16'hffdf;
  rom[20889] = 16'hffff;
  rom[20890] = 16'hffff;
  rom[20891] = 16'hffff;
  rom[20892] = 16'hf7bf;
  rom[20893] = 16'hf79f;
  rom[20894] = 16'hffff;
  rom[20895] = 16'hffff;
  rom[20896] = 16'hffff;
  rom[20897] = 16'hffff;
  rom[20898] = 16'hffff;
  rom[20899] = 16'hffff;
  rom[20900] = 16'hffdf;
  rom[20901] = 16'hffdf;
  rom[20902] = 16'hffff;
  rom[20903] = 16'hffff;
  rom[20904] = 16'hffff;
  rom[20905] = 16'hffff;
  rom[20906] = 16'hffff;
  rom[20907] = 16'hffff;
  rom[20908] = 16'hffff;
  rom[20909] = 16'hffff;
  rom[20910] = 16'hffff;
  rom[20911] = 16'hffff;
  rom[20912] = 16'hffff;
  rom[20913] = 16'hffff;
  rom[20914] = 16'hffff;
  rom[20915] = 16'hffff;
  rom[20916] = 16'hffff;
  rom[20917] = 16'hffff;
  rom[20918] = 16'hffff;
  rom[20919] = 16'hffff;
  rom[20920] = 16'hffff;
  rom[20921] = 16'hffff;
  rom[20922] = 16'hffff;
  rom[20923] = 16'hffff;
  rom[20924] = 16'hffff;
  rom[20925] = 16'hffff;
  rom[20926] = 16'hffff;
  rom[20927] = 16'hd656;
  rom[20928] = 16'h8b67;
  rom[20929] = 16'he54d;
  rom[20930] = 16'hf529;
  rom[20931] = 16'hfd48;
  rom[20932] = 16'hf506;
  rom[20933] = 16'hfd28;
  rom[20934] = 16'hfd08;
  rom[20935] = 16'hfd29;
  rom[20936] = 16'hfd08;
  rom[20937] = 16'hf509;
  rom[20938] = 16'hf528;
  rom[20939] = 16'hf54a;
  rom[20940] = 16'hf52a;
  rom[20941] = 16'hed2b;
  rom[20942] = 16'hdd0b;
  rom[20943] = 16'h82c4;
  rom[20944] = 16'h9c4c;
  rom[20945] = 16'hf73b;
  rom[20946] = 16'hffff;
  rom[20947] = 16'hffdf;
  rom[20948] = 16'hffff;
  rom[20949] = 16'hffff;
  rom[20950] = 16'hffff;
  rom[20951] = 16'hffff;
  rom[20952] = 16'hffff;
  rom[20953] = 16'hffff;
  rom[20954] = 16'hffff;
  rom[20955] = 16'hffff;
  rom[20956] = 16'hffff;
  rom[20957] = 16'hffff;
  rom[20958] = 16'hffff;
  rom[20959] = 16'hffff;
  rom[20960] = 16'hffff;
  rom[20961] = 16'hffff;
  rom[20962] = 16'hffff;
  rom[20963] = 16'hffff;
  rom[20964] = 16'hffff;
  rom[20965] = 16'hffff;
  rom[20966] = 16'hffff;
  rom[20967] = 16'hffff;
  rom[20968] = 16'hffff;
  rom[20969] = 16'hffff;
  rom[20970] = 16'hffff;
  rom[20971] = 16'hffff;
  rom[20972] = 16'hffff;
  rom[20973] = 16'hffff;
  rom[20974] = 16'hffff;
  rom[20975] = 16'hffff;
  rom[20976] = 16'hffff;
  rom[20977] = 16'hffff;
  rom[20978] = 16'hffff;
  rom[20979] = 16'hffff;
  rom[20980] = 16'hffff;
  rom[20981] = 16'hffff;
  rom[20982] = 16'hffff;
  rom[20983] = 16'hffff;
  rom[20984] = 16'hffff;
  rom[20985] = 16'hffff;
  rom[20986] = 16'hffff;
  rom[20987] = 16'hffff;
  rom[20988] = 16'hffff;
  rom[20989] = 16'hffff;
  rom[20990] = 16'hffff;
  rom[20991] = 16'hffff;
  rom[20992] = 16'hffff;
  rom[20993] = 16'hffff;
  rom[20994] = 16'hffff;
  rom[20995] = 16'hffff;
  rom[20996] = 16'hffff;
  rom[20997] = 16'hffff;
  rom[20998] = 16'hffff;
  rom[20999] = 16'hffff;
  rom[21000] = 16'hffff;
  rom[21001] = 16'hffff;
  rom[21002] = 16'hffff;
  rom[21003] = 16'hffff;
  rom[21004] = 16'hffff;
  rom[21005] = 16'hffff;
  rom[21006] = 16'hffff;
  rom[21007] = 16'hffff;
  rom[21008] = 16'hffff;
  rom[21009] = 16'hffff;
  rom[21010] = 16'hffff;
  rom[21011] = 16'hffff;
  rom[21012] = 16'hffff;
  rom[21013] = 16'hffff;
  rom[21014] = 16'hffff;
  rom[21015] = 16'hffff;
  rom[21016] = 16'hffff;
  rom[21017] = 16'hffff;
  rom[21018] = 16'hffff;
  rom[21019] = 16'hffff;
  rom[21020] = 16'hffff;
  rom[21021] = 16'hffff;
  rom[21022] = 16'hffff;
  rom[21023] = 16'hffff;
  rom[21024] = 16'hffff;
  rom[21025] = 16'hffff;
  rom[21026] = 16'hffff;
  rom[21027] = 16'hffff;
  rom[21028] = 16'hffff;
  rom[21029] = 16'hffff;
  rom[21030] = 16'hffff;
  rom[21031] = 16'hffff;
  rom[21032] = 16'hffff;
  rom[21033] = 16'hfffd;
  rom[21034] = 16'h9cad;
  rom[21035] = 16'h6b04;
  rom[21036] = 16'he68f;
  rom[21037] = 16'he6cb;
  rom[21038] = 16'hff8d;
  rom[21039] = 16'hf729;
  rom[21040] = 16'hff48;
  rom[21041] = 16'hf748;
  rom[21042] = 16'hf729;
  rom[21043] = 16'hf749;
  rom[21044] = 16'hf74a;
  rom[21045] = 16'hff29;
  rom[21046] = 16'hff2a;
  rom[21047] = 16'hff29;
  rom[21048] = 16'hff2a;
  rom[21049] = 16'hf729;
  rom[21050] = 16'hf74a;
  rom[21051] = 16'hef08;
  rom[21052] = 16'hff6a;
  rom[21053] = 16'hf70b;
  rom[21054] = 16'hee2c;
  rom[21055] = 16'h7a60;
  rom[21056] = 16'hab65;
  rom[21057] = 16'hed4c;
  rom[21058] = 16'hf529;
  rom[21059] = 16'hf507;
  rom[21060] = 16'hfd29;
  rom[21061] = 16'hfd09;
  rom[21062] = 16'hfd09;
  rom[21063] = 16'hfd69;
  rom[21064] = 16'he508;
  rom[21065] = 16'hd50a;
  rom[21066] = 16'h9ba9;
  rom[21067] = 16'hffde;
  rom[21068] = 16'hffff;
  rom[21069] = 16'hffff;
  rom[21070] = 16'hffff;
  rom[21071] = 16'hffff;
  rom[21072] = 16'hffff;
  rom[21073] = 16'hffff;
  rom[21074] = 16'hffff;
  rom[21075] = 16'hffff;
  rom[21076] = 16'hffff;
  rom[21077] = 16'hffff;
  rom[21078] = 16'hffff;
  rom[21079] = 16'hffff;
  rom[21080] = 16'hffff;
  rom[21081] = 16'hffff;
  rom[21082] = 16'hffff;
  rom[21083] = 16'hffff;
  rom[21084] = 16'hffff;
  rom[21085] = 16'hffff;
  rom[21086] = 16'hffff;
  rom[21087] = 16'hffff;
  rom[21088] = 16'hffff;
  rom[21089] = 16'hffff;
  rom[21090] = 16'hffff;
  rom[21091] = 16'hffff;
  rom[21092] = 16'hffff;
  rom[21093] = 16'hffff;
  rom[21094] = 16'hffff;
  rom[21095] = 16'hffff;
  rom[21096] = 16'hffff;
  rom[21097] = 16'hffff;
  rom[21098] = 16'hffff;
  rom[21099] = 16'hffff;
  rom[21100] = 16'hffff;
  rom[21101] = 16'hffff;
  rom[21102] = 16'hffff;
  rom[21103] = 16'hffff;
  rom[21104] = 16'hffff;
  rom[21105] = 16'hffff;
  rom[21106] = 16'hffff;
  rom[21107] = 16'hffff;
  rom[21108] = 16'hffff;
  rom[21109] = 16'hffff;
  rom[21110] = 16'hffff;
  rom[21111] = 16'hffff;
  rom[21112] = 16'hffff;
  rom[21113] = 16'hffff;
  rom[21114] = 16'hffff;
  rom[21115] = 16'hffff;
  rom[21116] = 16'hffff;
  rom[21117] = 16'hffff;
  rom[21118] = 16'hffff;
  rom[21119] = 16'hffff;
  rom[21120] = 16'hffff;
  rom[21121] = 16'hffff;
  rom[21122] = 16'hffff;
  rom[21123] = 16'hffff;
  rom[21124] = 16'hffff;
  rom[21125] = 16'hffff;
  rom[21126] = 16'hffde;
  rom[21127] = 16'hc5d3;
  rom[21128] = 16'h9ba9;
  rom[21129] = 16'he52c;
  rom[21130] = 16'hf50a;
  rom[21131] = 16'hfd07;
  rom[21132] = 16'hfd48;
  rom[21133] = 16'hfd07;
  rom[21134] = 16'hfd29;
  rom[21135] = 16'hfd09;
  rom[21136] = 16'hf508;
  rom[21137] = 16'hf528;
  rom[21138] = 16'hf4c8;
  rom[21139] = 16'hfd6b;
  rom[21140] = 16'hf54c;
  rom[21141] = 16'hd4cb;
  rom[21142] = 16'h9347;
  rom[21143] = 16'h8baa;
  rom[21144] = 16'hef39;
  rom[21145] = 16'hffff;
  rom[21146] = 16'hffff;
  rom[21147] = 16'hffff;
  rom[21148] = 16'hffff;
  rom[21149] = 16'hffff;
  rom[21150] = 16'hffff;
  rom[21151] = 16'hffff;
  rom[21152] = 16'hffff;
  rom[21153] = 16'hffff;
  rom[21154] = 16'hffff;
  rom[21155] = 16'hffff;
  rom[21156] = 16'hffff;
  rom[21157] = 16'hffff;
  rom[21158] = 16'hffff;
  rom[21159] = 16'hffff;
  rom[21160] = 16'hffff;
  rom[21161] = 16'hffff;
  rom[21162] = 16'hffff;
  rom[21163] = 16'hffff;
  rom[21164] = 16'hffff;
  rom[21165] = 16'hffff;
  rom[21166] = 16'hffff;
  rom[21167] = 16'hffff;
  rom[21168] = 16'hffff;
  rom[21169] = 16'hffff;
  rom[21170] = 16'hffff;
  rom[21171] = 16'hffff;
  rom[21172] = 16'hffff;
  rom[21173] = 16'hffff;
  rom[21174] = 16'hffff;
  rom[21175] = 16'hffff;
  rom[21176] = 16'hffff;
  rom[21177] = 16'hffff;
  rom[21178] = 16'hffff;
  rom[21179] = 16'hffff;
  rom[21180] = 16'hffff;
  rom[21181] = 16'hffff;
  rom[21182] = 16'hffff;
  rom[21183] = 16'hffff;
  rom[21184] = 16'hffff;
  rom[21185] = 16'hffff;
  rom[21186] = 16'hffff;
  rom[21187] = 16'hffff;
  rom[21188] = 16'hffff;
  rom[21189] = 16'hffff;
  rom[21190] = 16'hffff;
  rom[21191] = 16'hffff;
  rom[21192] = 16'hffff;
  rom[21193] = 16'hffff;
  rom[21194] = 16'hffff;
  rom[21195] = 16'hffff;
  rom[21196] = 16'hffff;
  rom[21197] = 16'hffff;
  rom[21198] = 16'hffff;
  rom[21199] = 16'hffff;
  rom[21200] = 16'hffff;
  rom[21201] = 16'hffff;
  rom[21202] = 16'hffff;
  rom[21203] = 16'hffff;
  rom[21204] = 16'hffff;
  rom[21205] = 16'hffff;
  rom[21206] = 16'hffff;
  rom[21207] = 16'hffff;
  rom[21208] = 16'hffff;
  rom[21209] = 16'hffff;
  rom[21210] = 16'hffff;
  rom[21211] = 16'hffff;
  rom[21212] = 16'hffff;
  rom[21213] = 16'hffff;
  rom[21214] = 16'hffff;
  rom[21215] = 16'hffff;
  rom[21216] = 16'hffff;
  rom[21217] = 16'hffff;
  rom[21218] = 16'hffff;
  rom[21219] = 16'hffff;
  rom[21220] = 16'hffff;
  rom[21221] = 16'hffff;
  rom[21222] = 16'hffff;
  rom[21223] = 16'hffff;
  rom[21224] = 16'hffff;
  rom[21225] = 16'hffff;
  rom[21226] = 16'hffff;
  rom[21227] = 16'hffff;
  rom[21228] = 16'hffff;
  rom[21229] = 16'hffff;
  rom[21230] = 16'hffff;
  rom[21231] = 16'hffff;
  rom[21232] = 16'hffde;
  rom[21233] = 16'hfffe;
  rom[21234] = 16'he739;
  rom[21235] = 16'h7b8a;
  rom[21236] = 16'h6ae5;
  rom[21237] = 16'heeaf;
  rom[21238] = 16'he6c9;
  rom[21239] = 16'hff48;
  rom[21240] = 16'hf727;
  rom[21241] = 16'hf729;
  rom[21242] = 16'hf729;
  rom[21243] = 16'hf72a;
  rom[21244] = 16'hf70a;
  rom[21245] = 16'hff0b;
  rom[21246] = 16'hf70a;
  rom[21247] = 16'hff29;
  rom[21248] = 16'hff09;
  rom[21249] = 16'hff29;
  rom[21250] = 16'hef29;
  rom[21251] = 16'hf749;
  rom[21252] = 16'hf748;
  rom[21253] = 16'hf6e9;
  rom[21254] = 16'hf6cb;
  rom[21255] = 16'hcd28;
  rom[21256] = 16'h7a61;
  rom[21257] = 16'hd4aa;
  rom[21258] = 16'hed48;
  rom[21259] = 16'hf547;
  rom[21260] = 16'hfd27;
  rom[21261] = 16'hfd2a;
  rom[21262] = 16'hf4c8;
  rom[21263] = 16'hfd28;
  rom[21264] = 16'hf548;
  rom[21265] = 16'hdd0b;
  rom[21266] = 16'h7265;
  rom[21267] = 16'hff7d;
  rom[21268] = 16'hffdf;
  rom[21269] = 16'hffff;
  rom[21270] = 16'hffff;
  rom[21271] = 16'hffff;
  rom[21272] = 16'hffff;
  rom[21273] = 16'hffff;
  rom[21274] = 16'hffff;
  rom[21275] = 16'hffff;
  rom[21276] = 16'hffff;
  rom[21277] = 16'hffff;
  rom[21278] = 16'hffff;
  rom[21279] = 16'hffff;
  rom[21280] = 16'hffff;
  rom[21281] = 16'hffff;
  rom[21282] = 16'hffff;
  rom[21283] = 16'hffff;
  rom[21284] = 16'hffff;
  rom[21285] = 16'hffff;
  rom[21286] = 16'hffff;
  rom[21287] = 16'hffff;
  rom[21288] = 16'hffff;
  rom[21289] = 16'hffff;
  rom[21290] = 16'hffff;
  rom[21291] = 16'hffff;
  rom[21292] = 16'hffff;
  rom[21293] = 16'hffff;
  rom[21294] = 16'hffff;
  rom[21295] = 16'hffff;
  rom[21296] = 16'hffff;
  rom[21297] = 16'hffff;
  rom[21298] = 16'hffff;
  rom[21299] = 16'hffff;
  rom[21300] = 16'hffff;
  rom[21301] = 16'hffff;
  rom[21302] = 16'hffff;
  rom[21303] = 16'hffff;
  rom[21304] = 16'hffff;
  rom[21305] = 16'hffff;
  rom[21306] = 16'hffff;
  rom[21307] = 16'hffff;
  rom[21308] = 16'hffff;
  rom[21309] = 16'hffff;
  rom[21310] = 16'hf7ff;
  rom[21311] = 16'hffff;
  rom[21312] = 16'hffff;
  rom[21313] = 16'hffff;
  rom[21314] = 16'hffff;
  rom[21315] = 16'hffff;
  rom[21316] = 16'hffff;
  rom[21317] = 16'hffff;
  rom[21318] = 16'hffff;
  rom[21319] = 16'hffff;
  rom[21320] = 16'hffff;
  rom[21321] = 16'hffff;
  rom[21322] = 16'hffff;
  rom[21323] = 16'hffff;
  rom[21324] = 16'hffff;
  rom[21325] = 16'hffff;
  rom[21326] = 16'hfffd;
  rom[21327] = 16'hb510;
  rom[21328] = 16'h9ba8;
  rom[21329] = 16'he54d;
  rom[21330] = 16'hf54a;
  rom[21331] = 16'hfd08;
  rom[21332] = 16'hfd07;
  rom[21333] = 16'hfd28;
  rom[21334] = 16'hfd08;
  rom[21335] = 16'hfd28;
  rom[21336] = 16'hfd28;
  rom[21337] = 16'hfd08;
  rom[21338] = 16'hf529;
  rom[21339] = 16'hed0b;
  rom[21340] = 16'hcc8a;
  rom[21341] = 16'h8b07;
  rom[21342] = 16'ha44d;
  rom[21343] = 16'hff7b;
  rom[21344] = 16'hfffe;
  rom[21345] = 16'hffff;
  rom[21346] = 16'hffff;
  rom[21347] = 16'hffff;
  rom[21348] = 16'hffff;
  rom[21349] = 16'hffff;
  rom[21350] = 16'hffff;
  rom[21351] = 16'hffff;
  rom[21352] = 16'hffff;
  rom[21353] = 16'hffff;
  rom[21354] = 16'hffff;
  rom[21355] = 16'hffff;
  rom[21356] = 16'hffff;
  rom[21357] = 16'hffff;
  rom[21358] = 16'hffff;
  rom[21359] = 16'hffff;
  rom[21360] = 16'hffff;
  rom[21361] = 16'hffff;
  rom[21362] = 16'hffff;
  rom[21363] = 16'hffff;
  rom[21364] = 16'hffff;
  rom[21365] = 16'hffff;
  rom[21366] = 16'hffff;
  rom[21367] = 16'hffff;
  rom[21368] = 16'hffff;
  rom[21369] = 16'hffff;
  rom[21370] = 16'hffff;
  rom[21371] = 16'hffff;
  rom[21372] = 16'hffff;
  rom[21373] = 16'hffff;
  rom[21374] = 16'hffff;
  rom[21375] = 16'hffff;
  rom[21376] = 16'hffff;
  rom[21377] = 16'hffff;
  rom[21378] = 16'hffff;
  rom[21379] = 16'hffff;
  rom[21380] = 16'hffff;
  rom[21381] = 16'hffff;
  rom[21382] = 16'hffff;
  rom[21383] = 16'hffff;
  rom[21384] = 16'hffff;
  rom[21385] = 16'hffff;
  rom[21386] = 16'hffff;
  rom[21387] = 16'hffff;
  rom[21388] = 16'hffff;
  rom[21389] = 16'hffff;
  rom[21390] = 16'hffff;
  rom[21391] = 16'hffff;
  rom[21392] = 16'hffff;
  rom[21393] = 16'hffff;
  rom[21394] = 16'hffff;
  rom[21395] = 16'hffff;
  rom[21396] = 16'hffff;
  rom[21397] = 16'hffff;
  rom[21398] = 16'hffff;
  rom[21399] = 16'hffff;
  rom[21400] = 16'hffff;
  rom[21401] = 16'hffff;
  rom[21402] = 16'hffff;
  rom[21403] = 16'hffff;
  rom[21404] = 16'hffff;
  rom[21405] = 16'hffff;
  rom[21406] = 16'hffff;
  rom[21407] = 16'hffff;
  rom[21408] = 16'hffff;
  rom[21409] = 16'hffff;
  rom[21410] = 16'hffff;
  rom[21411] = 16'hffff;
  rom[21412] = 16'hffff;
  rom[21413] = 16'hffff;
  rom[21414] = 16'hffff;
  rom[21415] = 16'hffff;
  rom[21416] = 16'hffff;
  rom[21417] = 16'hffff;
  rom[21418] = 16'hffff;
  rom[21419] = 16'hffff;
  rom[21420] = 16'hffff;
  rom[21421] = 16'hffff;
  rom[21422] = 16'hffff;
  rom[21423] = 16'hffff;
  rom[21424] = 16'hffff;
  rom[21425] = 16'hffff;
  rom[21426] = 16'hffff;
  rom[21427] = 16'hffff;
  rom[21428] = 16'hffff;
  rom[21429] = 16'hffff;
  rom[21430] = 16'hffff;
  rom[21431] = 16'hffff;
  rom[21432] = 16'hffff;
  rom[21433] = 16'hffff;
  rom[21434] = 16'hfffe;
  rom[21435] = 16'hdeda;
  rom[21436] = 16'h7329;
  rom[21437] = 16'h7b65;
  rom[21438] = 16'hf70d;
  rom[21439] = 16'hf769;
  rom[21440] = 16'hff48;
  rom[21441] = 16'hff28;
  rom[21442] = 16'hff2a;
  rom[21443] = 16'hf6c9;
  rom[21444] = 16'hff2b;
  rom[21445] = 16'hf70a;
  rom[21446] = 16'hff2a;
  rom[21447] = 16'hff29;
  rom[21448] = 16'hff2a;
  rom[21449] = 16'hf729;
  rom[21450] = 16'hff4a;
  rom[21451] = 16'hf727;
  rom[21452] = 16'hf727;
  rom[21453] = 16'hffaa;
  rom[21454] = 16'hf6ca;
  rom[21455] = 16'hf6ad;
  rom[21456] = 16'h9365;
  rom[21457] = 16'h82a0;
  rom[21458] = 16'he54a;
  rom[21459] = 16'hed48;
  rom[21460] = 16'hf508;
  rom[21461] = 16'hfd08;
  rom[21462] = 16'hfd08;
  rom[21463] = 16'hfd07;
  rom[21464] = 16'hfd49;
  rom[21465] = 16'hdcea;
  rom[21466] = 16'h7aa6;
  rom[21467] = 16'he659;
  rom[21468] = 16'hffff;
  rom[21469] = 16'hffff;
  rom[21470] = 16'hffff;
  rom[21471] = 16'hffff;
  rom[21472] = 16'hffff;
  rom[21473] = 16'hffff;
  rom[21474] = 16'hffff;
  rom[21475] = 16'hffff;
  rom[21476] = 16'hffff;
  rom[21477] = 16'hffff;
  rom[21478] = 16'hffff;
  rom[21479] = 16'hffff;
  rom[21480] = 16'hffff;
  rom[21481] = 16'hffff;
  rom[21482] = 16'hffff;
  rom[21483] = 16'hffff;
  rom[21484] = 16'hffff;
  rom[21485] = 16'hffff;
  rom[21486] = 16'hffff;
  rom[21487] = 16'hffff;
  rom[21488] = 16'hffff;
  rom[21489] = 16'hffff;
  rom[21490] = 16'hffff;
  rom[21491] = 16'hffff;
  rom[21492] = 16'hffff;
  rom[21493] = 16'hffff;
  rom[21494] = 16'hffff;
  rom[21495] = 16'hffff;
  rom[21496] = 16'hffff;
  rom[21497] = 16'hffff;
  rom[21498] = 16'hffff;
  rom[21499] = 16'hffff;
  rom[21500] = 16'hffff;
  rom[21501] = 16'hffff;
  rom[21502] = 16'hffff;
  rom[21503] = 16'hffff;
  rom[21504] = 16'hffff;
  rom[21505] = 16'hffff;
  rom[21506] = 16'hffff;
  rom[21507] = 16'hffff;
  rom[21508] = 16'hffff;
  rom[21509] = 16'hffff;
  rom[21510] = 16'hffff;
  rom[21511] = 16'hffff;
  rom[21512] = 16'hffff;
  rom[21513] = 16'hffff;
  rom[21514] = 16'hffff;
  rom[21515] = 16'hffff;
  rom[21516] = 16'hffff;
  rom[21517] = 16'hffff;
  rom[21518] = 16'hffff;
  rom[21519] = 16'hffff;
  rom[21520] = 16'hffff;
  rom[21521] = 16'hffff;
  rom[21522] = 16'hffff;
  rom[21523] = 16'hffff;
  rom[21524] = 16'hffff;
  rom[21525] = 16'hffff;
  rom[21526] = 16'hffdd;
  rom[21527] = 16'ha42c;
  rom[21528] = 16'hb46b;
  rom[21529] = 16'hed6d;
  rom[21530] = 16'hf52a;
  rom[21531] = 16'hfd07;
  rom[21532] = 16'hfd48;
  rom[21533] = 16'hfd07;
  rom[21534] = 16'hfd69;
  rom[21535] = 16'hf528;
  rom[21536] = 16'hfd29;
  rom[21537] = 16'hf52a;
  rom[21538] = 16'hed2b;
  rom[21539] = 16'hbc29;
  rom[21540] = 16'h6a03;
  rom[21541] = 16'haccf;
  rom[21542] = 16'hff9d;
  rom[21543] = 16'hffff;
  rom[21544] = 16'hffff;
  rom[21545] = 16'hffff;
  rom[21546] = 16'hffff;
  rom[21547] = 16'hffff;
  rom[21548] = 16'hffff;
  rom[21549] = 16'hffff;
  rom[21550] = 16'hffff;
  rom[21551] = 16'hffff;
  rom[21552] = 16'hffff;
  rom[21553] = 16'hffff;
  rom[21554] = 16'hffff;
  rom[21555] = 16'hffff;
  rom[21556] = 16'hffff;
  rom[21557] = 16'hffff;
  rom[21558] = 16'hffff;
  rom[21559] = 16'hffff;
  rom[21560] = 16'hffff;
  rom[21561] = 16'hffff;
  rom[21562] = 16'hffff;
  rom[21563] = 16'hffff;
  rom[21564] = 16'hffff;
  rom[21565] = 16'hffff;
  rom[21566] = 16'hffff;
  rom[21567] = 16'hffff;
  rom[21568] = 16'hffff;
  rom[21569] = 16'hffff;
  rom[21570] = 16'hffff;
  rom[21571] = 16'hffff;
  rom[21572] = 16'hffff;
  rom[21573] = 16'hffff;
  rom[21574] = 16'hffff;
  rom[21575] = 16'hffff;
  rom[21576] = 16'hffff;
  rom[21577] = 16'hffff;
  rom[21578] = 16'hffff;
  rom[21579] = 16'hffff;
  rom[21580] = 16'hffff;
  rom[21581] = 16'hffff;
  rom[21582] = 16'hffff;
  rom[21583] = 16'hffff;
  rom[21584] = 16'hffff;
  rom[21585] = 16'hffff;
  rom[21586] = 16'hffff;
  rom[21587] = 16'hffff;
  rom[21588] = 16'hffff;
  rom[21589] = 16'hffff;
  rom[21590] = 16'hffff;
  rom[21591] = 16'hffff;
  rom[21592] = 16'hffff;
  rom[21593] = 16'hffff;
  rom[21594] = 16'hffff;
  rom[21595] = 16'hffff;
  rom[21596] = 16'hffff;
  rom[21597] = 16'hffff;
  rom[21598] = 16'hffff;
  rom[21599] = 16'hffff;
  rom[21600] = 16'hffff;
  rom[21601] = 16'hffff;
  rom[21602] = 16'hffff;
  rom[21603] = 16'hffff;
  rom[21604] = 16'hffff;
  rom[21605] = 16'hffff;
  rom[21606] = 16'hffff;
  rom[21607] = 16'hffff;
  rom[21608] = 16'hffff;
  rom[21609] = 16'hffff;
  rom[21610] = 16'hffff;
  rom[21611] = 16'hffff;
  rom[21612] = 16'hffff;
  rom[21613] = 16'hffff;
  rom[21614] = 16'hffff;
  rom[21615] = 16'hffff;
  rom[21616] = 16'hffff;
  rom[21617] = 16'hffff;
  rom[21618] = 16'hffff;
  rom[21619] = 16'hffff;
  rom[21620] = 16'hffff;
  rom[21621] = 16'hffff;
  rom[21622] = 16'hffff;
  rom[21623] = 16'hffff;
  rom[21624] = 16'hffff;
  rom[21625] = 16'hffff;
  rom[21626] = 16'hffff;
  rom[21627] = 16'hffff;
  rom[21628] = 16'hffff;
  rom[21629] = 16'hffff;
  rom[21630] = 16'hffff;
  rom[21631] = 16'hffff;
  rom[21632] = 16'hffff;
  rom[21633] = 16'hffff;
  rom[21634] = 16'hffff;
  rom[21635] = 16'hffff;
  rom[21636] = 16'he6da;
  rom[21637] = 16'h62a6;
  rom[21638] = 16'h8be5;
  rom[21639] = 16'heeab;
  rom[21640] = 16'hf729;
  rom[21641] = 16'hff29;
  rom[21642] = 16'hff09;
  rom[21643] = 16'hff2a;
  rom[21644] = 16'hff09;
  rom[21645] = 16'hff29;
  rom[21646] = 16'hf729;
  rom[21647] = 16'hff29;
  rom[21648] = 16'hf729;
  rom[21649] = 16'hf729;
  rom[21650] = 16'hf729;
  rom[21651] = 16'hf748;
  rom[21652] = 16'hef47;
  rom[21653] = 16'hf749;
  rom[21654] = 16'hf72a;
  rom[21655] = 16'hfeed;
  rom[21656] = 16'hcd69;
  rom[21657] = 16'h7280;
  rom[21658] = 16'ha3a4;
  rom[21659] = 16'hf56a;
  rom[21660] = 16'hf529;
  rom[21661] = 16'hfd08;
  rom[21662] = 16'hfd07;
  rom[21663] = 16'hfd07;
  rom[21664] = 16'hf4e7;
  rom[21665] = 16'hed4c;
  rom[21666] = 16'ha3c9;
  rom[21667] = 16'h9c4e;
  rom[21668] = 16'hffbd;
  rom[21669] = 16'hffff;
  rom[21670] = 16'hffff;
  rom[21671] = 16'hffff;
  rom[21672] = 16'hffff;
  rom[21673] = 16'hffff;
  rom[21674] = 16'hffff;
  rom[21675] = 16'hffff;
  rom[21676] = 16'hffff;
  rom[21677] = 16'hffff;
  rom[21678] = 16'hffff;
  rom[21679] = 16'hffff;
  rom[21680] = 16'hffff;
  rom[21681] = 16'hffff;
  rom[21682] = 16'hffdf;
  rom[21683] = 16'hffff;
  rom[21684] = 16'hffff;
  rom[21685] = 16'hffff;
  rom[21686] = 16'hf7ff;
  rom[21687] = 16'hffff;
  rom[21688] = 16'hffff;
  rom[21689] = 16'hffff;
  rom[21690] = 16'hffff;
  rom[21691] = 16'hffff;
  rom[21692] = 16'hffdf;
  rom[21693] = 16'hffff;
  rom[21694] = 16'hffff;
  rom[21695] = 16'hffff;
  rom[21696] = 16'hffde;
  rom[21697] = 16'hffff;
  rom[21698] = 16'hffff;
  rom[21699] = 16'hffff;
  rom[21700] = 16'hffff;
  rom[21701] = 16'hffff;
  rom[21702] = 16'hffff;
  rom[21703] = 16'hffff;
  rom[21704] = 16'hffff;
  rom[21705] = 16'hffff;
  rom[21706] = 16'hffff;
  rom[21707] = 16'hffff;
  rom[21708] = 16'hffff;
  rom[21709] = 16'hffff;
  rom[21710] = 16'hffff;
  rom[21711] = 16'hffff;
  rom[21712] = 16'hffdf;
  rom[21713] = 16'hffff;
  rom[21714] = 16'hffff;
  rom[21715] = 16'hffff;
  rom[21716] = 16'hffff;
  rom[21717] = 16'hffff;
  rom[21718] = 16'hffff;
  rom[21719] = 16'hffff;
  rom[21720] = 16'hffff;
  rom[21721] = 16'hffff;
  rom[21722] = 16'hffff;
  rom[21723] = 16'hffff;
  rom[21724] = 16'hffff;
  rom[21725] = 16'hffff;
  rom[21726] = 16'hf6fa;
  rom[21727] = 16'h8308;
  rom[21728] = 16'hc4ab;
  rom[21729] = 16'hed2b;
  rom[21730] = 16'hf528;
  rom[21731] = 16'hfd47;
  rom[21732] = 16'hf527;
  rom[21733] = 16'hf548;
  rom[21734] = 16'hed28;
  rom[21735] = 16'hed6a;
  rom[21736] = 16'hed6c;
  rom[21737] = 16'hd4cb;
  rom[21738] = 16'ha3a7;
  rom[21739] = 16'h8b28;
  rom[21740] = 16'hbd93;
  rom[21741] = 16'hffde;
  rom[21742] = 16'hffbf;
  rom[21743] = 16'hffff;
  rom[21744] = 16'hffdf;
  rom[21745] = 16'hffdf;
  rom[21746] = 16'hffff;
  rom[21747] = 16'hffff;
  rom[21748] = 16'hffff;
  rom[21749] = 16'hffff;
  rom[21750] = 16'hffff;
  rom[21751] = 16'hffff;
  rom[21752] = 16'hffff;
  rom[21753] = 16'hffff;
  rom[21754] = 16'hffff;
  rom[21755] = 16'hffff;
  rom[21756] = 16'hffff;
  rom[21757] = 16'hffff;
  rom[21758] = 16'hffff;
  rom[21759] = 16'hffff;
  rom[21760] = 16'hffff;
  rom[21761] = 16'hffff;
  rom[21762] = 16'hffff;
  rom[21763] = 16'hffff;
  rom[21764] = 16'hffff;
  rom[21765] = 16'hffff;
  rom[21766] = 16'hffff;
  rom[21767] = 16'hffff;
  rom[21768] = 16'hffff;
  rom[21769] = 16'hffff;
  rom[21770] = 16'hffff;
  rom[21771] = 16'hffff;
  rom[21772] = 16'hffff;
  rom[21773] = 16'hffff;
  rom[21774] = 16'hffff;
  rom[21775] = 16'hffff;
  rom[21776] = 16'hffff;
  rom[21777] = 16'hffff;
  rom[21778] = 16'hffff;
  rom[21779] = 16'hffff;
  rom[21780] = 16'hffff;
  rom[21781] = 16'hffff;
  rom[21782] = 16'hffff;
  rom[21783] = 16'hffff;
  rom[21784] = 16'hffff;
  rom[21785] = 16'hffff;
  rom[21786] = 16'hffff;
  rom[21787] = 16'hffff;
  rom[21788] = 16'hffff;
  rom[21789] = 16'hffff;
  rom[21790] = 16'hffff;
  rom[21791] = 16'hffff;
  rom[21792] = 16'hffff;
  rom[21793] = 16'hffff;
  rom[21794] = 16'hffff;
  rom[21795] = 16'hffff;
  rom[21796] = 16'hffff;
  rom[21797] = 16'hffff;
  rom[21798] = 16'hffff;
  rom[21799] = 16'hffff;
  rom[21800] = 16'hffff;
  rom[21801] = 16'hffff;
  rom[21802] = 16'hffff;
  rom[21803] = 16'hffff;
  rom[21804] = 16'hffff;
  rom[21805] = 16'hffff;
  rom[21806] = 16'hffff;
  rom[21807] = 16'hffff;
  rom[21808] = 16'hffff;
  rom[21809] = 16'hffff;
  rom[21810] = 16'hffff;
  rom[21811] = 16'hffff;
  rom[21812] = 16'hffff;
  rom[21813] = 16'hffff;
  rom[21814] = 16'hffff;
  rom[21815] = 16'hffff;
  rom[21816] = 16'hffff;
  rom[21817] = 16'hffff;
  rom[21818] = 16'hffff;
  rom[21819] = 16'hffff;
  rom[21820] = 16'hffff;
  rom[21821] = 16'hffff;
  rom[21822] = 16'hffff;
  rom[21823] = 16'hffff;
  rom[21824] = 16'hffff;
  rom[21825] = 16'hffff;
  rom[21826] = 16'hffff;
  rom[21827] = 16'hffff;
  rom[21828] = 16'hffff;
  rom[21829] = 16'hffff;
  rom[21830] = 16'hffff;
  rom[21831] = 16'hffff;
  rom[21832] = 16'hffff;
  rom[21833] = 16'hffff;
  rom[21834] = 16'hffff;
  rom[21835] = 16'hffff;
  rom[21836] = 16'hffdf;
  rom[21837] = 16'hde98;
  rom[21838] = 16'h41c3;
  rom[21839] = 16'h83a5;
  rom[21840] = 16'he66c;
  rom[21841] = 16'hf70c;
  rom[21842] = 16'hfeea;
  rom[21843] = 16'hff4a;
  rom[21844] = 16'hff28;
  rom[21845] = 16'hff48;
  rom[21846] = 16'hff49;
  rom[21847] = 16'hf728;
  rom[21848] = 16'hff49;
  rom[21849] = 16'hf728;
  rom[21850] = 16'hff49;
  rom[21851] = 16'hf728;
  rom[21852] = 16'hef07;
  rom[21853] = 16'hf729;
  rom[21854] = 16'hf72b;
  rom[21855] = 16'hf6eb;
  rom[21856] = 16'hf6cd;
  rom[21857] = 16'hb4e7;
  rom[21858] = 16'h7a62;
  rom[21859] = 16'hcc69;
  rom[21860] = 16'hf54b;
  rom[21861] = 16'hf529;
  rom[21862] = 16'hf4a5;
  rom[21863] = 16'hfd07;
  rom[21864] = 16'hfd2a;
  rom[21865] = 16'hed2c;
  rom[21866] = 16'hc4ab;
  rom[21867] = 16'h6aa5;
  rom[21868] = 16'hef1a;
  rom[21869] = 16'hffff;
  rom[21870] = 16'hffff;
  rom[21871] = 16'hffbf;
  rom[21872] = 16'hffff;
  rom[21873] = 16'hffff;
  rom[21874] = 16'hffff;
  rom[21875] = 16'hffff;
  rom[21876] = 16'hffff;
  rom[21877] = 16'hffff;
  rom[21878] = 16'hffff;
  rom[21879] = 16'hffff;
  rom[21880] = 16'hffff;
  rom[21881] = 16'hffff;
  rom[21882] = 16'hffff;
  rom[21883] = 16'hffff;
  rom[21884] = 16'hffff;
  rom[21885] = 16'hffff;
  rom[21886] = 16'hffff;
  rom[21887] = 16'hffff;
  rom[21888] = 16'hffff;
  rom[21889] = 16'hffdf;
  rom[21890] = 16'hffbf;
  rom[21891] = 16'hffbe;
  rom[21892] = 16'hffff;
  rom[21893] = 16'hffff;
  rom[21894] = 16'hffff;
  rom[21895] = 16'hffff;
  rom[21896] = 16'hffff;
  rom[21897] = 16'hffff;
  rom[21898] = 16'hffff;
  rom[21899] = 16'hffff;
  rom[21900] = 16'hffff;
  rom[21901] = 16'hfffe;
  rom[21902] = 16'hffff;
  rom[21903] = 16'hffde;
  rom[21904] = 16'hffff;
  rom[21905] = 16'hffff;
  rom[21906] = 16'hffdf;
  rom[21907] = 16'hffdf;
  rom[21908] = 16'hffdf;
  rom[21909] = 16'hffdf;
  rom[21910] = 16'hffdf;
  rom[21911] = 16'hffdf;
  rom[21912] = 16'hffff;
  rom[21913] = 16'hffff;
  rom[21914] = 16'hffff;
  rom[21915] = 16'hffff;
  rom[21916] = 16'hffff;
  rom[21917] = 16'hffff;
  rom[21918] = 16'hffff;
  rom[21919] = 16'hffff;
  rom[21920] = 16'hffff;
  rom[21921] = 16'hffff;
  rom[21922] = 16'hffff;
  rom[21923] = 16'hffff;
  rom[21924] = 16'hffff;
  rom[21925] = 16'hffff;
  rom[21926] = 16'hac70;
  rom[21927] = 16'h9b48;
  rom[21928] = 16'hdcec;
  rom[21929] = 16'he529;
  rom[21930] = 16'hfd89;
  rom[21931] = 16'hf527;
  rom[21932] = 16'hfd28;
  rom[21933] = 16'he507;
  rom[21934] = 16'hed6b;
  rom[21935] = 16'hdd6c;
  rom[21936] = 16'hc4ab;
  rom[21937] = 16'h82c6;
  rom[21938] = 16'h93ab;
  rom[21939] = 16'he6d8;
  rom[21940] = 16'hffde;
  rom[21941] = 16'hf7df;
  rom[21942] = 16'hffff;
  rom[21943] = 16'hffff;
  rom[21944] = 16'hffff;
  rom[21945] = 16'hffff;
  rom[21946] = 16'hffff;
  rom[21947] = 16'hffff;
  rom[21948] = 16'hffff;
  rom[21949] = 16'hffff;
  rom[21950] = 16'hffff;
  rom[21951] = 16'hffff;
  rom[21952] = 16'hffff;
  rom[21953] = 16'hffff;
  rom[21954] = 16'hffff;
  rom[21955] = 16'hffff;
  rom[21956] = 16'hffff;
  rom[21957] = 16'hffff;
  rom[21958] = 16'hffff;
  rom[21959] = 16'hffff;
  rom[21960] = 16'hffff;
  rom[21961] = 16'hffff;
  rom[21962] = 16'hffff;
  rom[21963] = 16'hffff;
  rom[21964] = 16'hffff;
  rom[21965] = 16'hffff;
  rom[21966] = 16'hffff;
  rom[21967] = 16'hffff;
  rom[21968] = 16'hffff;
  rom[21969] = 16'hffff;
  rom[21970] = 16'hffff;
  rom[21971] = 16'hffff;
  rom[21972] = 16'hffff;
  rom[21973] = 16'hffff;
  rom[21974] = 16'hffff;
  rom[21975] = 16'hffff;
  rom[21976] = 16'hffff;
  rom[21977] = 16'hffff;
  rom[21978] = 16'hffff;
  rom[21979] = 16'hffff;
  rom[21980] = 16'hffff;
  rom[21981] = 16'hffff;
  rom[21982] = 16'hffff;
  rom[21983] = 16'hffff;
  rom[21984] = 16'hffff;
  rom[21985] = 16'hffff;
  rom[21986] = 16'hffff;
  rom[21987] = 16'hffff;
  rom[21988] = 16'hffff;
  rom[21989] = 16'hffff;
  rom[21990] = 16'hffff;
  rom[21991] = 16'hffff;
  rom[21992] = 16'hffff;
  rom[21993] = 16'hffff;
  rom[21994] = 16'hffff;
  rom[21995] = 16'hffff;
  rom[21996] = 16'hffff;
  rom[21997] = 16'hffff;
  rom[21998] = 16'hffff;
  rom[21999] = 16'hffff;
  rom[22000] = 16'hffff;
  rom[22001] = 16'hffff;
  rom[22002] = 16'hffff;
  rom[22003] = 16'hffff;
  rom[22004] = 16'hffff;
  rom[22005] = 16'hffff;
  rom[22006] = 16'hffff;
  rom[22007] = 16'hffff;
  rom[22008] = 16'hffff;
  rom[22009] = 16'hffff;
  rom[22010] = 16'hffff;
  rom[22011] = 16'hffff;
  rom[22012] = 16'hffff;
  rom[22013] = 16'hffff;
  rom[22014] = 16'hffff;
  rom[22015] = 16'hffff;
  rom[22016] = 16'hffff;
  rom[22017] = 16'hffff;
  rom[22018] = 16'hffff;
  rom[22019] = 16'hffff;
  rom[22020] = 16'hffff;
  rom[22021] = 16'hffff;
  rom[22022] = 16'hffff;
  rom[22023] = 16'hffff;
  rom[22024] = 16'hffff;
  rom[22025] = 16'hffff;
  rom[22026] = 16'hffff;
  rom[22027] = 16'hffff;
  rom[22028] = 16'hffff;
  rom[22029] = 16'hffff;
  rom[22030] = 16'hffff;
  rom[22031] = 16'hffff;
  rom[22032] = 16'hffff;
  rom[22033] = 16'hffff;
  rom[22034] = 16'hffff;
  rom[22035] = 16'hffff;
  rom[22036] = 16'hffff;
  rom[22037] = 16'hffff;
  rom[22038] = 16'he6fa;
  rom[22039] = 16'h5a65;
  rom[22040] = 16'h8c07;
  rom[22041] = 16'hde2d;
  rom[22042] = 16'hf74e;
  rom[22043] = 16'heec8;
  rom[22044] = 16'hf748;
  rom[22045] = 16'hff69;
  rom[22046] = 16'hf707;
  rom[22047] = 16'hff49;
  rom[22048] = 16'hf708;
  rom[22049] = 16'hff49;
  rom[22050] = 16'hef28;
  rom[22051] = 16'hf728;
  rom[22052] = 16'hff29;
  rom[22053] = 16'hff4a;
  rom[22054] = 16'hef09;
  rom[22055] = 16'hff2b;
  rom[22056] = 16'hf72c;
  rom[22057] = 16'hf6ac;
  rom[22058] = 16'h93a4;
  rom[22059] = 16'h7a61;
  rom[22060] = 16'hcceb;
  rom[22061] = 16'he52a;
  rom[22062] = 16'hfdcb;
  rom[22063] = 16'hfd09;
  rom[22064] = 16'hfcea;
  rom[22065] = 16'hf56d;
  rom[22066] = 16'hdd4c;
  rom[22067] = 16'h7b04;
  rom[22068] = 16'hc573;
  rom[22069] = 16'hfffe;
  rom[22070] = 16'hffde;
  rom[22071] = 16'hffff;
  rom[22072] = 16'hffff;
  rom[22073] = 16'hffff;
  rom[22074] = 16'hffff;
  rom[22075] = 16'hffff;
  rom[22076] = 16'hffff;
  rom[22077] = 16'hffff;
  rom[22078] = 16'hffff;
  rom[22079] = 16'hffff;
  rom[22080] = 16'hffff;
  rom[22081] = 16'hffff;
  rom[22082] = 16'hffff;
  rom[22083] = 16'hffff;
  rom[22084] = 16'hffff;
  rom[22085] = 16'hffff;
  rom[22086] = 16'hffff;
  rom[22087] = 16'hffff;
  rom[22088] = 16'hff9d;
  rom[22089] = 16'hf6bb;
  rom[22090] = 16'hff3c;
  rom[22091] = 16'hff9d;
  rom[22092] = 16'hffdd;
  rom[22093] = 16'hffde;
  rom[22094] = 16'hffbd;
  rom[22095] = 16'hffde;
  rom[22096] = 16'hfffe;
  rom[22097] = 16'hfffe;
  rom[22098] = 16'hffde;
  rom[22099] = 16'hffde;
  rom[22100] = 16'hffbd;
  rom[22101] = 16'hffde;
  rom[22102] = 16'hff9c;
  rom[22103] = 16'hff3c;
  rom[22104] = 16'hf6fa;
  rom[22105] = 16'heedb;
  rom[22106] = 16'hffdf;
  rom[22107] = 16'hffff;
  rom[22108] = 16'hffdf;
  rom[22109] = 16'hffff;
  rom[22110] = 16'hffdf;
  rom[22111] = 16'hffff;
  rom[22112] = 16'hffff;
  rom[22113] = 16'hffff;
  rom[22114] = 16'hffff;
  rom[22115] = 16'hffff;
  rom[22116] = 16'hffff;
  rom[22117] = 16'hffff;
  rom[22118] = 16'hffff;
  rom[22119] = 16'hffff;
  rom[22120] = 16'hffff;
  rom[22121] = 16'hffff;
  rom[22122] = 16'hffff;
  rom[22123] = 16'hffff;
  rom[22124] = 16'hffff;
  rom[22125] = 16'hf73c;
  rom[22126] = 16'h8b29;
  rom[22127] = 16'hbc2b;
  rom[22128] = 16'he50b;
  rom[22129] = 16'hf56a;
  rom[22130] = 16'hf508;
  rom[22131] = 16'hfd49;
  rom[22132] = 16'hf529;
  rom[22133] = 16'hf5ad;
  rom[22134] = 16'hc4ca;
  rom[22135] = 16'h9ba9;
  rom[22136] = 16'h7ae8;
  rom[22137] = 16'hbd33;
  rom[22138] = 16'hffde;
  rom[22139] = 16'hffff;
  rom[22140] = 16'hffff;
  rom[22141] = 16'hffff;
  rom[22142] = 16'hffff;
  rom[22143] = 16'hffff;
  rom[22144] = 16'hffff;
  rom[22145] = 16'hffff;
  rom[22146] = 16'hffff;
  rom[22147] = 16'hffff;
  rom[22148] = 16'hffff;
  rom[22149] = 16'hffff;
  rom[22150] = 16'hffff;
  rom[22151] = 16'hffff;
  rom[22152] = 16'hffff;
  rom[22153] = 16'hffff;
  rom[22154] = 16'hffff;
  rom[22155] = 16'hffff;
  rom[22156] = 16'hffff;
  rom[22157] = 16'hffff;
  rom[22158] = 16'hffff;
  rom[22159] = 16'hffff;
  rom[22160] = 16'hffff;
  rom[22161] = 16'hffff;
  rom[22162] = 16'hffff;
  rom[22163] = 16'hffff;
  rom[22164] = 16'hffff;
  rom[22165] = 16'hffff;
  rom[22166] = 16'hffff;
  rom[22167] = 16'hffff;
  rom[22168] = 16'hffff;
  rom[22169] = 16'hffff;
  rom[22170] = 16'hffff;
  rom[22171] = 16'hffff;
  rom[22172] = 16'hffff;
  rom[22173] = 16'hffff;
  rom[22174] = 16'hffff;
  rom[22175] = 16'hffff;
  rom[22176] = 16'hffff;
  rom[22177] = 16'hffff;
  rom[22178] = 16'hffff;
  rom[22179] = 16'hffff;
  rom[22180] = 16'hffff;
  rom[22181] = 16'hffff;
  rom[22182] = 16'hffff;
  rom[22183] = 16'hffff;
  rom[22184] = 16'hffff;
  rom[22185] = 16'hffff;
  rom[22186] = 16'hffff;
  rom[22187] = 16'hffff;
  rom[22188] = 16'hffff;
  rom[22189] = 16'hffff;
  rom[22190] = 16'hffff;
  rom[22191] = 16'hffff;
  rom[22192] = 16'hffff;
  rom[22193] = 16'hffff;
  rom[22194] = 16'hffff;
  rom[22195] = 16'hffff;
  rom[22196] = 16'hffff;
  rom[22197] = 16'hffff;
  rom[22198] = 16'hffff;
  rom[22199] = 16'hffff;
  rom[22200] = 16'hffff;
  rom[22201] = 16'hffff;
  rom[22202] = 16'hffff;
  rom[22203] = 16'hffff;
  rom[22204] = 16'hffff;
  rom[22205] = 16'hffff;
  rom[22206] = 16'hffff;
  rom[22207] = 16'hffff;
  rom[22208] = 16'hffff;
  rom[22209] = 16'hffff;
  rom[22210] = 16'hffff;
  rom[22211] = 16'hffff;
  rom[22212] = 16'hffff;
  rom[22213] = 16'hffff;
  rom[22214] = 16'hffff;
  rom[22215] = 16'hffff;
  rom[22216] = 16'hffff;
  rom[22217] = 16'hffff;
  rom[22218] = 16'hffff;
  rom[22219] = 16'hffff;
  rom[22220] = 16'hffff;
  rom[22221] = 16'hffff;
  rom[22222] = 16'hffff;
  rom[22223] = 16'hffff;
  rom[22224] = 16'hffff;
  rom[22225] = 16'hffff;
  rom[22226] = 16'hffff;
  rom[22227] = 16'hffff;
  rom[22228] = 16'hffff;
  rom[22229] = 16'hffff;
  rom[22230] = 16'hffff;
  rom[22231] = 16'hffff;
  rom[22232] = 16'hffff;
  rom[22233] = 16'hffff;
  rom[22234] = 16'hffff;
  rom[22235] = 16'hffff;
  rom[22236] = 16'hffdf;
  rom[22237] = 16'hffff;
  rom[22238] = 16'hffff;
  rom[22239] = 16'hd697;
  rom[22240] = 16'h7328;
  rom[22241] = 16'h7b66;
  rom[22242] = 16'hd60c;
  rom[22243] = 16'hf74d;
  rom[22244] = 16'hef29;
  rom[22245] = 16'hf748;
  rom[22246] = 16'hff49;
  rom[22247] = 16'hf729;
  rom[22248] = 16'hff4a;
  rom[22249] = 16'hf728;
  rom[22250] = 16'hf749;
  rom[22251] = 16'hf728;
  rom[22252] = 16'hff29;
  rom[22253] = 16'hf709;
  rom[22254] = 16'hff4a;
  rom[22255] = 16'hef08;
  rom[22256] = 16'hf729;
  rom[22257] = 16'hff4b;
  rom[22258] = 16'hde0b;
  rom[22259] = 16'h7ae2;
  rom[22260] = 16'h82c4;
  rom[22261] = 16'hc4aa;
  rom[22262] = 16'hdceb;
  rom[22263] = 16'hed2b;
  rom[22264] = 16'hfd2c;
  rom[22265] = 16'he4ea;
  rom[22266] = 16'hdd2c;
  rom[22267] = 16'hbccc;
  rom[22268] = 16'h836a;
  rom[22269] = 16'hffbd;
  rom[22270] = 16'hffff;
  rom[22271] = 16'hffff;
  rom[22272] = 16'hffff;
  rom[22273] = 16'hffff;
  rom[22274] = 16'hffff;
  rom[22275] = 16'hffff;
  rom[22276] = 16'hffff;
  rom[22277] = 16'hffff;
  rom[22278] = 16'hffff;
  rom[22279] = 16'hffff;
  rom[22280] = 16'hffff;
  rom[22281] = 16'hffff;
  rom[22282] = 16'hffff;
  rom[22283] = 16'hffff;
  rom[22284] = 16'hffff;
  rom[22285] = 16'hffff;
  rom[22286] = 16'hffff;
  rom[22287] = 16'hffde;
  rom[22288] = 16'hff7e;
  rom[22289] = 16'hc4d3;
  rom[22290] = 16'hc450;
  rom[22291] = 16'hdcf2;
  rom[22292] = 16'hf5b5;
  rom[22293] = 16'hfe17;
  rom[22294] = 16'hfed9;
  rom[22295] = 16'hfef9;
  rom[22296] = 16'hff1b;
  rom[22297] = 16'hfed9;
  rom[22298] = 16'hff1a;
  rom[22299] = 16'hfefa;
  rom[22300] = 16'hfe78;
  rom[22301] = 16'hedb6;
  rom[22302] = 16'he554;
  rom[22303] = 16'hcc71;
  rom[22304] = 16'hbc50;
  rom[22305] = 16'hddd7;
  rom[22306] = 16'hffbe;
  rom[22307] = 16'hffdf;
  rom[22308] = 16'hffff;
  rom[22309] = 16'hffff;
  rom[22310] = 16'hffff;
  rom[22311] = 16'hffff;
  rom[22312] = 16'hffff;
  rom[22313] = 16'hffff;
  rom[22314] = 16'hffff;
  rom[22315] = 16'hffff;
  rom[22316] = 16'hffff;
  rom[22317] = 16'hffff;
  rom[22318] = 16'hffff;
  rom[22319] = 16'hffff;
  rom[22320] = 16'hffff;
  rom[22321] = 16'hffff;
  rom[22322] = 16'hffff;
  rom[22323] = 16'hffff;
  rom[22324] = 16'hfffe;
  rom[22325] = 16'hbd72;
  rom[22326] = 16'h8b07;
  rom[22327] = 16'hdcec;
  rom[22328] = 16'hed2b;
  rom[22329] = 16'hf528;
  rom[22330] = 16'hf508;
  rom[22331] = 16'hfd0a;
  rom[22332] = 16'heceb;
  rom[22333] = 16'hab88;
  rom[22334] = 16'h82c7;
  rom[22335] = 16'hb48f;
  rom[22336] = 16'he699;
  rom[22337] = 16'hff9f;
  rom[22338] = 16'hffff;
  rom[22339] = 16'hffff;
  rom[22340] = 16'hffff;
  rom[22341] = 16'hffff;
  rom[22342] = 16'hffff;
  rom[22343] = 16'hffff;
  rom[22344] = 16'hffff;
  rom[22345] = 16'hffff;
  rom[22346] = 16'hffff;
  rom[22347] = 16'hffff;
  rom[22348] = 16'hffff;
  rom[22349] = 16'hffff;
  rom[22350] = 16'hffff;
  rom[22351] = 16'hffff;
  rom[22352] = 16'hffff;
  rom[22353] = 16'hffff;
  rom[22354] = 16'hffff;
  rom[22355] = 16'hffff;
  rom[22356] = 16'hffff;
  rom[22357] = 16'hffff;
  rom[22358] = 16'hffff;
  rom[22359] = 16'hffff;
  rom[22360] = 16'hffff;
  rom[22361] = 16'hffff;
  rom[22362] = 16'hffff;
  rom[22363] = 16'hffff;
  rom[22364] = 16'hffff;
  rom[22365] = 16'hffff;
  rom[22366] = 16'hffff;
  rom[22367] = 16'hffff;
  rom[22368] = 16'hffff;
  rom[22369] = 16'hffff;
  rom[22370] = 16'hffff;
  rom[22371] = 16'hffff;
  rom[22372] = 16'hffff;
  rom[22373] = 16'hffff;
  rom[22374] = 16'hffff;
  rom[22375] = 16'hffff;
  rom[22376] = 16'hffff;
  rom[22377] = 16'hffff;
  rom[22378] = 16'hffff;
  rom[22379] = 16'hffff;
  rom[22380] = 16'hffff;
  rom[22381] = 16'hffff;
  rom[22382] = 16'hffff;
  rom[22383] = 16'hffff;
  rom[22384] = 16'hffff;
  rom[22385] = 16'hffff;
  rom[22386] = 16'hffff;
  rom[22387] = 16'hffff;
  rom[22388] = 16'hffff;
  rom[22389] = 16'hffff;
  rom[22390] = 16'hffff;
  rom[22391] = 16'hffff;
  rom[22392] = 16'hffff;
  rom[22393] = 16'hffff;
  rom[22394] = 16'hffff;
  rom[22395] = 16'hffff;
  rom[22396] = 16'hffff;
  rom[22397] = 16'hffff;
  rom[22398] = 16'hffff;
  rom[22399] = 16'hffff;
  rom[22400] = 16'hffff;
  rom[22401] = 16'hffff;
  rom[22402] = 16'hffff;
  rom[22403] = 16'hffff;
  rom[22404] = 16'hffff;
  rom[22405] = 16'hffff;
  rom[22406] = 16'hffff;
  rom[22407] = 16'hffff;
  rom[22408] = 16'hffff;
  rom[22409] = 16'hffff;
  rom[22410] = 16'hffff;
  rom[22411] = 16'hffff;
  rom[22412] = 16'hffff;
  rom[22413] = 16'hffff;
  rom[22414] = 16'hffff;
  rom[22415] = 16'hffff;
  rom[22416] = 16'hffff;
  rom[22417] = 16'hffff;
  rom[22418] = 16'hffff;
  rom[22419] = 16'hffff;
  rom[22420] = 16'hffff;
  rom[22421] = 16'hffff;
  rom[22422] = 16'hffff;
  rom[22423] = 16'hffff;
  rom[22424] = 16'hffff;
  rom[22425] = 16'hffff;
  rom[22426] = 16'hffff;
  rom[22427] = 16'hffff;
  rom[22428] = 16'hffff;
  rom[22429] = 16'hffff;
  rom[22430] = 16'hffff;
  rom[22431] = 16'hffff;
  rom[22432] = 16'hffff;
  rom[22433] = 16'hffff;
  rom[22434] = 16'hffff;
  rom[22435] = 16'hffff;
  rom[22436] = 16'hffde;
  rom[22437] = 16'hffff;
  rom[22438] = 16'hffff;
  rom[22439] = 16'hfffe;
  rom[22440] = 16'hf79b;
  rom[22441] = 16'h62e7;
  rom[22442] = 16'h6b24;
  rom[22443] = 16'hc5ea;
  rom[22444] = 16'hef2c;
  rom[22445] = 16'hef0a;
  rom[22446] = 16'hff4a;
  rom[22447] = 16'hf70a;
  rom[22448] = 16'hf729;
  rom[22449] = 16'hff29;
  rom[22450] = 16'hff08;
  rom[22451] = 16'hff09;
  rom[22452] = 16'hf709;
  rom[22453] = 16'hf729;
  rom[22454] = 16'hf728;
  rom[22455] = 16'hff88;
  rom[22456] = 16'hef27;
  rom[22457] = 16'hf6e8;
  rom[22458] = 16'hf6ec;
  rom[22459] = 16'hcdcb;
  rom[22460] = 16'h6241;
  rom[22461] = 16'h61e2;
  rom[22462] = 16'ha347;
  rom[22463] = 16'hc3c8;
  rom[22464] = 16'hdc6a;
  rom[22465] = 16'hf54d;
  rom[22466] = 16'he52d;
  rom[22467] = 16'hdd90;
  rom[22468] = 16'h7b08;
  rom[22469] = 16'ha490;
  rom[22470] = 16'hffbe;
  rom[22471] = 16'hffff;
  rom[22472] = 16'hffff;
  rom[22473] = 16'hffff;
  rom[22474] = 16'hffff;
  rom[22475] = 16'hffff;
  rom[22476] = 16'hffff;
  rom[22477] = 16'hffff;
  rom[22478] = 16'hffff;
  rom[22479] = 16'hffff;
  rom[22480] = 16'hffff;
  rom[22481] = 16'hffff;
  rom[22482] = 16'hffff;
  rom[22483] = 16'hffff;
  rom[22484] = 16'hffff;
  rom[22485] = 16'hffff;
  rom[22486] = 16'hffdf;
  rom[22487] = 16'hffff;
  rom[22488] = 16'hffbd;
  rom[22489] = 16'hedf7;
  rom[22490] = 16'hab0b;
  rom[22491] = 16'hbaca;
  rom[22492] = 16'hbaea;
  rom[22493] = 16'hc2e9;
  rom[22494] = 16'hbac9;
  rom[22495] = 16'hbaa9;
  rom[22496] = 16'hbac9;
  rom[22497] = 16'hc2e9;
  rom[22498] = 16'hb2c8;
  rom[22499] = 16'hc2e9;
  rom[22500] = 16'hc30a;
  rom[22501] = 16'hc2ea;
  rom[22502] = 16'hbaca;
  rom[22503] = 16'hb2eb;
  rom[22504] = 16'hcc50;
  rom[22505] = 16'hff7d;
  rom[22506] = 16'hffde;
  rom[22507] = 16'hffff;
  rom[22508] = 16'hffff;
  rom[22509] = 16'hffff;
  rom[22510] = 16'hffff;
  rom[22511] = 16'hffff;
  rom[22512] = 16'hffff;
  rom[22513] = 16'hffff;
  rom[22514] = 16'hffff;
  rom[22515] = 16'hffff;
  rom[22516] = 16'hffff;
  rom[22517] = 16'hffff;
  rom[22518] = 16'hffff;
  rom[22519] = 16'hffff;
  rom[22520] = 16'hffff;
  rom[22521] = 16'hffff;
  rom[22522] = 16'hffdf;
  rom[22523] = 16'hffff;
  rom[22524] = 16'hd697;
  rom[22525] = 16'h8baa;
  rom[22526] = 16'hbc6b;
  rom[22527] = 16'hed0b;
  rom[22528] = 16'hece9;
  rom[22529] = 16'hfd09;
  rom[22530] = 16'heca8;
  rom[22531] = 16'hcba6;
  rom[22532] = 16'h8a02;
  rom[22533] = 16'h71e4;
  rom[22534] = 16'he5d5;
  rom[22535] = 16'hff3b;
  rom[22536] = 16'hffbd;
  rom[22537] = 16'hffbf;
  rom[22538] = 16'hff9e;
  rom[22539] = 16'hffdf;
  rom[22540] = 16'hfffe;
  rom[22541] = 16'hffdd;
  rom[22542] = 16'hfffe;
  rom[22543] = 16'hffff;
  rom[22544] = 16'hffde;
  rom[22545] = 16'hffff;
  rom[22546] = 16'hffff;
  rom[22547] = 16'hffff;
  rom[22548] = 16'hffff;
  rom[22549] = 16'hffff;
  rom[22550] = 16'hffff;
  rom[22551] = 16'hffff;
  rom[22552] = 16'hffff;
  rom[22553] = 16'hffff;
  rom[22554] = 16'hffff;
  rom[22555] = 16'hffff;
  rom[22556] = 16'hffff;
  rom[22557] = 16'hffff;
  rom[22558] = 16'hffff;
  rom[22559] = 16'hffff;
  rom[22560] = 16'hffff;
  rom[22561] = 16'hffff;
  rom[22562] = 16'hffff;
  rom[22563] = 16'hffff;
  rom[22564] = 16'hffff;
  rom[22565] = 16'hffff;
  rom[22566] = 16'hffff;
  rom[22567] = 16'hffff;
  rom[22568] = 16'hffff;
  rom[22569] = 16'hffff;
  rom[22570] = 16'hffff;
  rom[22571] = 16'hffff;
  rom[22572] = 16'hffff;
  rom[22573] = 16'hffff;
  rom[22574] = 16'hffff;
  rom[22575] = 16'hffff;
  rom[22576] = 16'hffff;
  rom[22577] = 16'hffff;
  rom[22578] = 16'hffff;
  rom[22579] = 16'hffff;
  rom[22580] = 16'hffff;
  rom[22581] = 16'hffff;
  rom[22582] = 16'hffff;
  rom[22583] = 16'hffff;
  rom[22584] = 16'hffff;
  rom[22585] = 16'hffff;
  rom[22586] = 16'hffff;
  rom[22587] = 16'hffff;
  rom[22588] = 16'hffff;
  rom[22589] = 16'hffff;
  rom[22590] = 16'hffff;
  rom[22591] = 16'hffff;
  rom[22592] = 16'hffff;
  rom[22593] = 16'hffff;
  rom[22594] = 16'hffff;
  rom[22595] = 16'hffff;
  rom[22596] = 16'hffff;
  rom[22597] = 16'hffff;
  rom[22598] = 16'hffff;
  rom[22599] = 16'hffff;
  rom[22600] = 16'hffff;
  rom[22601] = 16'hffff;
  rom[22602] = 16'hffff;
  rom[22603] = 16'hffff;
  rom[22604] = 16'hffff;
  rom[22605] = 16'hffff;
  rom[22606] = 16'hffff;
  rom[22607] = 16'hffff;
  rom[22608] = 16'hffff;
  rom[22609] = 16'hffff;
  rom[22610] = 16'hffff;
  rom[22611] = 16'hffff;
  rom[22612] = 16'hffff;
  rom[22613] = 16'hffff;
  rom[22614] = 16'hffff;
  rom[22615] = 16'hffff;
  rom[22616] = 16'hffff;
  rom[22617] = 16'hffff;
  rom[22618] = 16'hffff;
  rom[22619] = 16'hffff;
  rom[22620] = 16'hffff;
  rom[22621] = 16'hffff;
  rom[22622] = 16'hffff;
  rom[22623] = 16'hffff;
  rom[22624] = 16'hffff;
  rom[22625] = 16'hffff;
  rom[22626] = 16'hffff;
  rom[22627] = 16'hffff;
  rom[22628] = 16'hffff;
  rom[22629] = 16'hffff;
  rom[22630] = 16'hffff;
  rom[22631] = 16'hffff;
  rom[22632] = 16'hffff;
  rom[22633] = 16'hffff;
  rom[22634] = 16'hffff;
  rom[22635] = 16'hffdf;
  rom[22636] = 16'hffdf;
  rom[22637] = 16'hffdf;
  rom[22638] = 16'hffff;
  rom[22639] = 16'hffff;
  rom[22640] = 16'hffff;
  rom[22641] = 16'he73b;
  rom[22642] = 16'h944d;
  rom[22643] = 16'h62c4;
  rom[22644] = 16'hb509;
  rom[22645] = 16'he6cd;
  rom[22646] = 16'hf70d;
  rom[22647] = 16'hf70b;
  rom[22648] = 16'hff2a;
  rom[22649] = 16'hfee9;
  rom[22650] = 16'hff0a;
  rom[22651] = 16'hff0a;
  rom[22652] = 16'hff4b;
  rom[22653] = 16'hef29;
  rom[22654] = 16'hf748;
  rom[22655] = 16'hf727;
  rom[22656] = 16'hff68;
  rom[22657] = 16'hf729;
  rom[22658] = 16'hff2b;
  rom[22659] = 16'hf72e;
  rom[22660] = 16'hcdab;
  rom[22661] = 16'h7282;
  rom[22662] = 16'h6160;
  rom[22663] = 16'h9244;
  rom[22664] = 16'h9243;
  rom[22665] = 16'h9aa4;
  rom[22666] = 16'hc3ca;
  rom[22667] = 16'hbbea;
  rom[22668] = 16'hb42c;
  rom[22669] = 16'h6266;
  rom[22670] = 16'hd5f7;
  rom[22671] = 16'hffdf;
  rom[22672] = 16'hffff;
  rom[22673] = 16'hffff;
  rom[22674] = 16'hffff;
  rom[22675] = 16'hffff;
  rom[22676] = 16'hffff;
  rom[22677] = 16'hffff;
  rom[22678] = 16'hffff;
  rom[22679] = 16'hffff;
  rom[22680] = 16'hffff;
  rom[22681] = 16'hffff;
  rom[22682] = 16'hffff;
  rom[22683] = 16'hffff;
  rom[22684] = 16'hffff;
  rom[22685] = 16'hffff;
  rom[22686] = 16'hffff;
  rom[22687] = 16'hffdf;
  rom[22688] = 16'hfffe;
  rom[22689] = 16'hff5c;
  rom[22690] = 16'hf595;
  rom[22691] = 16'hcb8c;
  rom[22692] = 16'hcae9;
  rom[22693] = 16'hca86;
  rom[22694] = 16'he2a8;
  rom[22695] = 16'hda66;
  rom[22696] = 16'hda87;
  rom[22697] = 16'hda87;
  rom[22698] = 16'hda88;
  rom[22699] = 16'hdaa8;
  rom[22700] = 16'hdaa9;
  rom[22701] = 16'hcaa8;
  rom[22702] = 16'hcaea;
  rom[22703] = 16'he491;
  rom[22704] = 16'hfeb9;
  rom[22705] = 16'hffbd;
  rom[22706] = 16'hfffe;
  rom[22707] = 16'hffff;
  rom[22708] = 16'hffff;
  rom[22709] = 16'hffff;
  rom[22710] = 16'hffff;
  rom[22711] = 16'hffff;
  rom[22712] = 16'hffff;
  rom[22713] = 16'hffff;
  rom[22714] = 16'hffff;
  rom[22715] = 16'hffff;
  rom[22716] = 16'hffff;
  rom[22717] = 16'hffff;
  rom[22718] = 16'hffff;
  rom[22719] = 16'hffff;
  rom[22720] = 16'hffff;
  rom[22721] = 16'hffff;
  rom[22722] = 16'hffdf;
  rom[22723] = 16'hf73d;
  rom[22724] = 16'h9c70;
  rom[22725] = 16'h8b6a;
  rom[22726] = 16'hed4f;
  rom[22727] = 16'hf4aa;
  rom[22728] = 16'hfc49;
  rom[22729] = 16'he366;
  rom[22730] = 16'hcb06;
  rom[22731] = 16'h9a23;
  rom[22732] = 16'h9ac5;
  rom[22733] = 16'h8265;
  rom[22734] = 16'h9b69;
  rom[22735] = 16'hb46d;
  rom[22736] = 16'hd5d4;
  rom[22737] = 16'he657;
  rom[22738] = 16'hf6fa;
  rom[22739] = 16'hff5c;
  rom[22740] = 16'hff9d;
  rom[22741] = 16'hffbe;
  rom[22742] = 16'hffdf;
  rom[22743] = 16'hffdf;
  rom[22744] = 16'hffff;
  rom[22745] = 16'hffff;
  rom[22746] = 16'hffff;
  rom[22747] = 16'hffff;
  rom[22748] = 16'hffff;
  rom[22749] = 16'hffff;
  rom[22750] = 16'hffff;
  rom[22751] = 16'hffff;
  rom[22752] = 16'hffff;
  rom[22753] = 16'hffff;
  rom[22754] = 16'hffff;
  rom[22755] = 16'hffff;
  rom[22756] = 16'hffff;
  rom[22757] = 16'hffff;
  rom[22758] = 16'hffff;
  rom[22759] = 16'hffff;
  rom[22760] = 16'hffff;
  rom[22761] = 16'hffff;
  rom[22762] = 16'hffff;
  rom[22763] = 16'hffff;
  rom[22764] = 16'hffff;
  rom[22765] = 16'hffff;
  rom[22766] = 16'hffff;
  rom[22767] = 16'hffff;
  rom[22768] = 16'hffff;
  rom[22769] = 16'hffff;
  rom[22770] = 16'hffff;
  rom[22771] = 16'hffff;
  rom[22772] = 16'hffff;
  rom[22773] = 16'hffff;
  rom[22774] = 16'hffff;
  rom[22775] = 16'hffff;
  rom[22776] = 16'hffff;
  rom[22777] = 16'hffff;
  rom[22778] = 16'hffff;
  rom[22779] = 16'hffff;
  rom[22780] = 16'hffff;
  rom[22781] = 16'hffff;
  rom[22782] = 16'hffff;
  rom[22783] = 16'hffff;
  rom[22784] = 16'hffff;
  rom[22785] = 16'hffff;
  rom[22786] = 16'hffff;
  rom[22787] = 16'hffff;
  rom[22788] = 16'hffff;
  rom[22789] = 16'hffff;
  rom[22790] = 16'hffff;
  rom[22791] = 16'hffff;
  rom[22792] = 16'hffff;
  rom[22793] = 16'hffff;
  rom[22794] = 16'hffff;
  rom[22795] = 16'hffff;
  rom[22796] = 16'hffff;
  rom[22797] = 16'hffff;
  rom[22798] = 16'hffff;
  rom[22799] = 16'hffff;
  rom[22800] = 16'hffff;
  rom[22801] = 16'hffff;
  rom[22802] = 16'hffff;
  rom[22803] = 16'hffff;
  rom[22804] = 16'hffff;
  rom[22805] = 16'hffff;
  rom[22806] = 16'hffff;
  rom[22807] = 16'hffff;
  rom[22808] = 16'hffff;
  rom[22809] = 16'hffff;
  rom[22810] = 16'hffff;
  rom[22811] = 16'hffff;
  rom[22812] = 16'hffff;
  rom[22813] = 16'hffff;
  rom[22814] = 16'hffff;
  rom[22815] = 16'hffff;
  rom[22816] = 16'hffff;
  rom[22817] = 16'hffff;
  rom[22818] = 16'hffff;
  rom[22819] = 16'hffff;
  rom[22820] = 16'hffff;
  rom[22821] = 16'hffff;
  rom[22822] = 16'hffff;
  rom[22823] = 16'hffff;
  rom[22824] = 16'hffff;
  rom[22825] = 16'hffff;
  rom[22826] = 16'hffff;
  rom[22827] = 16'hffff;
  rom[22828] = 16'hffff;
  rom[22829] = 16'hffff;
  rom[22830] = 16'hffff;
  rom[22831] = 16'hffff;
  rom[22832] = 16'hffff;
  rom[22833] = 16'hffff;
  rom[22834] = 16'hffff;
  rom[22835] = 16'hffff;
  rom[22836] = 16'hffbf;
  rom[22837] = 16'hffdf;
  rom[22838] = 16'hffde;
  rom[22839] = 16'hffff;
  rom[22840] = 16'hffff;
  rom[22841] = 16'hffff;
  rom[22842] = 16'hf7be;
  rom[22843] = 16'hbd92;
  rom[22844] = 16'h5aa4;
  rom[22845] = 16'h9406;
  rom[22846] = 16'heeee;
  rom[22847] = 16'hef0d;
  rom[22848] = 16'heeeb;
  rom[22849] = 16'hff4b;
  rom[22850] = 16'hfee9;
  rom[22851] = 16'hff09;
  rom[22852] = 16'hf708;
  rom[22853] = 16'hff8b;
  rom[22854] = 16'hef28;
  rom[22855] = 16'hf769;
  rom[22856] = 16'hf728;
  rom[22857] = 16'hff49;
  rom[22858] = 16'hef29;
  rom[22859] = 16'hef0a;
  rom[22860] = 16'hf72c;
  rom[22861] = 16'hddca;
  rom[22862] = 16'h8ac1;
  rom[22863] = 16'h9aa3;
  rom[22864] = 16'haae6;
  rom[22865] = 16'haaa6;
  rom[22866] = 16'h9a24;
  rom[22867] = 16'h8161;
  rom[22868] = 16'h8a04;
  rom[22869] = 16'h8247;
  rom[22870] = 16'h6227;
  rom[22871] = 16'hf6fb;
  rom[22872] = 16'hffbf;
  rom[22873] = 16'hffff;
  rom[22874] = 16'hffdf;
  rom[22875] = 16'hffff;
  rom[22876] = 16'hffdf;
  rom[22877] = 16'hffff;
  rom[22878] = 16'hffff;
  rom[22879] = 16'hffff;
  rom[22880] = 16'hffff;
  rom[22881] = 16'hffff;
  rom[22882] = 16'hffff;
  rom[22883] = 16'hffff;
  rom[22884] = 16'hffff;
  rom[22885] = 16'hffff;
  rom[22886] = 16'hffff;
  rom[22887] = 16'hfffe;
  rom[22888] = 16'hffde;
  rom[22889] = 16'hfffd;
  rom[22890] = 16'hff9a;
  rom[22891] = 16'hf5f4;
  rom[22892] = 16'hd40d;
  rom[22893] = 16'hc2c8;
  rom[22894] = 16'hd2a7;
  rom[22895] = 16'he287;
  rom[22896] = 16'he2a8;
  rom[22897] = 16'hda87;
  rom[22898] = 16'hd288;
  rom[22899] = 16'hd268;
  rom[22900] = 16'hd267;
  rom[22901] = 16'hd34b;
  rom[22902] = 16'hdc6f;
  rom[22903] = 16'hfed8;
  rom[22904] = 16'hffbc;
  rom[22905] = 16'hfffe;
  rom[22906] = 16'hf7fd;
  rom[22907] = 16'hf7fe;
  rom[22908] = 16'hffff;
  rom[22909] = 16'hffff;
  rom[22910] = 16'hffff;
  rom[22911] = 16'hffff;
  rom[22912] = 16'hffff;
  rom[22913] = 16'hffff;
  rom[22914] = 16'hffff;
  rom[22915] = 16'hffff;
  rom[22916] = 16'hffff;
  rom[22917] = 16'hffff;
  rom[22918] = 16'hffff;
  rom[22919] = 16'hffff;
  rom[22920] = 16'hffff;
  rom[22921] = 16'hffff;
  rom[22922] = 16'hff9d;
  rom[22923] = 16'hb4b2;
  rom[22924] = 16'h7a88;
  rom[22925] = 16'hc42d;
  rom[22926] = 16'hdbeb;
  rom[22927] = 16'hdb06;
  rom[22928] = 16'he2c5;
  rom[22929] = 16'hd283;
  rom[22930] = 16'hcac4;
  rom[22931] = 16'haae3;
  rom[22932] = 16'hc407;
  rom[22933] = 16'h92e3;
  rom[22934] = 16'h82c1;
  rom[22935] = 16'h6a41;
  rom[22936] = 16'h49c1;
  rom[22937] = 16'h6243;
  rom[22938] = 16'h6244;
  rom[22939] = 16'ha42c;
  rom[22940] = 16'hc511;
  rom[22941] = 16'he617;
  rom[22942] = 16'hfefa;
  rom[22943] = 16'hff5c;
  rom[22944] = 16'hff5d;
  rom[22945] = 16'hffdf;
  rom[22946] = 16'hffbe;
  rom[22947] = 16'hffde;
  rom[22948] = 16'hffff;
  rom[22949] = 16'hffff;
  rom[22950] = 16'hfffe;
  rom[22951] = 16'hffff;
  rom[22952] = 16'hffff;
  rom[22953] = 16'hffff;
  rom[22954] = 16'hffdf;
  rom[22955] = 16'hffff;
  rom[22956] = 16'hffff;
  rom[22957] = 16'hffff;
  rom[22958] = 16'hffff;
  rom[22959] = 16'hffff;
  rom[22960] = 16'hffff;
  rom[22961] = 16'hffff;
  rom[22962] = 16'hffff;
  rom[22963] = 16'hffff;
  rom[22964] = 16'hffff;
  rom[22965] = 16'hffff;
  rom[22966] = 16'hffff;
  rom[22967] = 16'hffff;
  rom[22968] = 16'hffff;
  rom[22969] = 16'hffff;
  rom[22970] = 16'hffff;
  rom[22971] = 16'hffff;
  rom[22972] = 16'hffff;
  rom[22973] = 16'hffff;
  rom[22974] = 16'hffdf;
  rom[22975] = 16'hffff;
  rom[22976] = 16'hffff;
  rom[22977] = 16'hffff;
  rom[22978] = 16'hffff;
  rom[22979] = 16'hffff;
  rom[22980] = 16'hffff;
  rom[22981] = 16'hffff;
  rom[22982] = 16'hffff;
  rom[22983] = 16'hffff;
  rom[22984] = 16'hffff;
  rom[22985] = 16'hffff;
  rom[22986] = 16'hffff;
  rom[22987] = 16'hffff;
  rom[22988] = 16'hffff;
  rom[22989] = 16'hffff;
  rom[22990] = 16'hffff;
  rom[22991] = 16'hffff;
  rom[22992] = 16'hffff;
  rom[22993] = 16'hffff;
  rom[22994] = 16'hffff;
  rom[22995] = 16'hffff;
  rom[22996] = 16'hffff;
  rom[22997] = 16'hffff;
  rom[22998] = 16'hffff;
  rom[22999] = 16'hffff;
  rom[23000] = 16'hffff;
  rom[23001] = 16'hffff;
  rom[23002] = 16'hffff;
  rom[23003] = 16'hffff;
  rom[23004] = 16'hffff;
  rom[23005] = 16'hffff;
  rom[23006] = 16'hffff;
  rom[23007] = 16'hffff;
  rom[23008] = 16'hffff;
  rom[23009] = 16'hffff;
  rom[23010] = 16'hffff;
  rom[23011] = 16'hffff;
  rom[23012] = 16'hffff;
  rom[23013] = 16'hffff;
  rom[23014] = 16'hffff;
  rom[23015] = 16'hffff;
  rom[23016] = 16'hffff;
  rom[23017] = 16'hffff;
  rom[23018] = 16'hffff;
  rom[23019] = 16'hffff;
  rom[23020] = 16'hffff;
  rom[23021] = 16'hffff;
  rom[23022] = 16'hffff;
  rom[23023] = 16'hffff;
  rom[23024] = 16'hffff;
  rom[23025] = 16'hffff;
  rom[23026] = 16'hffff;
  rom[23027] = 16'hffff;
  rom[23028] = 16'hffff;
  rom[23029] = 16'hffff;
  rom[23030] = 16'hffff;
  rom[23031] = 16'hffff;
  rom[23032] = 16'hffff;
  rom[23033] = 16'hffff;
  rom[23034] = 16'hffff;
  rom[23035] = 16'hffdf;
  rom[23036] = 16'hffdf;
  rom[23037] = 16'hffff;
  rom[23038] = 16'hffff;
  rom[23039] = 16'hffff;
  rom[23040] = 16'hffff;
  rom[23041] = 16'hffdf;
  rom[23042] = 16'hffff;
  rom[23043] = 16'hffde;
  rom[23044] = 16'hce14;
  rom[23045] = 16'h7346;
  rom[23046] = 16'h7b65;
  rom[23047] = 16'hc60c;
  rom[23048] = 16'hef2f;
  rom[23049] = 16'heeeb;
  rom[23050] = 16'hff6c;
  rom[23051] = 16'hf708;
  rom[23052] = 16'hff4a;
  rom[23053] = 16'hef08;
  rom[23054] = 16'hf749;
  rom[23055] = 16'hf709;
  rom[23056] = 16'hf729;
  rom[23057] = 16'hf729;
  rom[23058] = 16'hff29;
  rom[23059] = 16'hff69;
  rom[23060] = 16'hf709;
  rom[23061] = 16'hff2c;
  rom[23062] = 16'hf60b;
  rom[23063] = 16'hc466;
  rom[23064] = 16'hb325;
  rom[23065] = 16'hb2a5;
  rom[23066] = 16'hc2e7;
  rom[23067] = 16'hc2a7;
  rom[23068] = 16'hc2a8;
  rom[23069] = 16'h99e5;
  rom[23070] = 16'h79e6;
  rom[23071] = 16'h936d;
  rom[23072] = 16'he67a;
  rom[23073] = 16'hffdf;
  rom[23074] = 16'hffdf;
  rom[23075] = 16'hffff;
  rom[23076] = 16'hffff;
  rom[23077] = 16'hffff;
  rom[23078] = 16'hffdf;
  rom[23079] = 16'hffff;
  rom[23080] = 16'hffff;
  rom[23081] = 16'hffff;
  rom[23082] = 16'hffff;
  rom[23083] = 16'hffff;
  rom[23084] = 16'hffff;
  rom[23085] = 16'hffff;
  rom[23086] = 16'hffff;
  rom[23087] = 16'hffff;
  rom[23088] = 16'hffff;
  rom[23089] = 16'hffdd;
  rom[23090] = 16'hfffd;
  rom[23091] = 16'hffbc;
  rom[23092] = 16'hff19;
  rom[23093] = 16'hf593;
  rom[23094] = 16'he44e;
  rom[23095] = 16'hd38b;
  rom[23096] = 16'hd36b;
  rom[23097] = 16'hd36b;
  rom[23098] = 16'hd3ad;
  rom[23099] = 16'hdbee;
  rom[23100] = 16'hfcf2;
  rom[23101] = 16'hfe37;
  rom[23102] = 16'hff1a;
  rom[23103] = 16'hffdd;
  rom[23104] = 16'hfffe;
  rom[23105] = 16'hfffe;
  rom[23106] = 16'hffff;
  rom[23107] = 16'hffff;
  rom[23108] = 16'hffff;
  rom[23109] = 16'hffff;
  rom[23110] = 16'hffff;
  rom[23111] = 16'hffff;
  rom[23112] = 16'hffff;
  rom[23113] = 16'hffff;
  rom[23114] = 16'hffff;
  rom[23115] = 16'hffdf;
  rom[23116] = 16'hffff;
  rom[23117] = 16'hffdf;
  rom[23118] = 16'hffff;
  rom[23119] = 16'hf7be;
  rom[23120] = 16'hffff;
  rom[23121] = 16'hff7c;
  rom[23122] = 16'hd554;
  rom[23123] = 16'h8247;
  rom[23124] = 16'ha266;
  rom[23125] = 16'hcb28;
  rom[23126] = 16'hcae7;
  rom[23127] = 16'hd2a5;
  rom[23128] = 16'hdaa4;
  rom[23129] = 16'hcae3;
  rom[23130] = 16'hd3e5;
  rom[23131] = 16'hfe0c;
  rom[23132] = 16'hfe4c;
  rom[23133] = 16'hfead;
  rom[23134] = 16'hfead;
  rom[23135] = 16'hcda9;
  rom[23136] = 16'hbd69;
  rom[23137] = 16'h9c66;
  rom[23138] = 16'h8b85;
  rom[23139] = 16'h6a42;
  rom[23140] = 16'h7222;
  rom[23141] = 16'h7243;
  rom[23142] = 16'h8ac7;
  rom[23143] = 16'ha3ac;
  rom[23144] = 16'hc4d1;
  rom[23145] = 16'hd553;
  rom[23146] = 16'hedf7;
  rom[23147] = 16'hee38;
  rom[23148] = 16'hfeb9;
  rom[23149] = 16'hfefa;
  rom[23150] = 16'hff3c;
  rom[23151] = 16'hff5c;
  rom[23152] = 16'hff7e;
  rom[23153] = 16'hffbf;
  rom[23154] = 16'hffbf;
  rom[23155] = 16'hffbf;
  rom[23156] = 16'hffdf;
  rom[23157] = 16'hffde;
  rom[23158] = 16'hffdf;
  rom[23159] = 16'hffdf;
  rom[23160] = 16'hffff;
  rom[23161] = 16'hffff;
  rom[23162] = 16'hffff;
  rom[23163] = 16'hffdf;
  rom[23164] = 16'hffff;
  rom[23165] = 16'hffdf;
  rom[23166] = 16'hffff;
  rom[23167] = 16'hffde;
  rom[23168] = 16'hffff;
  rom[23169] = 16'hffff;
  rom[23170] = 16'hffbe;
  rom[23171] = 16'hffbe;
  rom[23172] = 16'hffbe;
  rom[23173] = 16'hff7d;
  rom[23174] = 16'hff1c;
  rom[23175] = 16'hfefb;
  rom[23176] = 16'hffbd;
  rom[23177] = 16'hffff;
  rom[23178] = 16'hffff;
  rom[23179] = 16'hffff;
  rom[23180] = 16'hffff;
  rom[23181] = 16'hffff;
  rom[23182] = 16'hffff;
  rom[23183] = 16'hffff;
  rom[23184] = 16'hffff;
  rom[23185] = 16'hffff;
  rom[23186] = 16'hffff;
  rom[23187] = 16'hffff;
  rom[23188] = 16'hffff;
  rom[23189] = 16'hffff;
  rom[23190] = 16'hffff;
  rom[23191] = 16'hffff;
  rom[23192] = 16'hffff;
  rom[23193] = 16'hffff;
  rom[23194] = 16'hffff;
  rom[23195] = 16'hffff;
  rom[23196] = 16'hffff;
  rom[23197] = 16'hffff;
  rom[23198] = 16'hffff;
  rom[23199] = 16'hffff;
  rom[23200] = 16'hffdf;
  rom[23201] = 16'hffff;
  rom[23202] = 16'hffff;
  rom[23203] = 16'hffff;
  rom[23204] = 16'hf7ff;
  rom[23205] = 16'hffff;
  rom[23206] = 16'hffff;
  rom[23207] = 16'hffff;
  rom[23208] = 16'hffff;
  rom[23209] = 16'hffff;
  rom[23210] = 16'hffdf;
  rom[23211] = 16'hffff;
  rom[23212] = 16'hffff;
  rom[23213] = 16'hffff;
  rom[23214] = 16'hffff;
  rom[23215] = 16'hffff;
  rom[23216] = 16'hf7ff;
  rom[23217] = 16'hffff;
  rom[23218] = 16'hffff;
  rom[23219] = 16'hffff;
  rom[23220] = 16'hffff;
  rom[23221] = 16'hffff;
  rom[23222] = 16'hffff;
  rom[23223] = 16'hffff;
  rom[23224] = 16'hffff;
  rom[23225] = 16'hffff;
  rom[23226] = 16'hffff;
  rom[23227] = 16'hffff;
  rom[23228] = 16'hffff;
  rom[23229] = 16'hffff;
  rom[23230] = 16'hffff;
  rom[23231] = 16'hffff;
  rom[23232] = 16'hffff;
  rom[23233] = 16'hffff;
  rom[23234] = 16'hffff;
  rom[23235] = 16'hffff;
  rom[23236] = 16'hffdf;
  rom[23237] = 16'hffff;
  rom[23238] = 16'hffff;
  rom[23239] = 16'hffff;
  rom[23240] = 16'hffdf;
  rom[23241] = 16'hffff;
  rom[23242] = 16'hffdf;
  rom[23243] = 16'hffdf;
  rom[23244] = 16'hffde;
  rom[23245] = 16'he6b9;
  rom[23246] = 16'h942c;
  rom[23247] = 16'h62e4;
  rom[23248] = 16'h9cc8;
  rom[23249] = 16'he6cd;
  rom[23250] = 16'he6ea;
  rom[23251] = 16'hff29;
  rom[23252] = 16'hf6e7;
  rom[23253] = 16'hff49;
  rom[23254] = 16'hf729;
  rom[23255] = 16'hff2a;
  rom[23256] = 16'hff29;
  rom[23257] = 16'hfee8;
  rom[23258] = 16'hf708;
  rom[23259] = 16'hff29;
  rom[23260] = 16'hf728;
  rom[23261] = 16'hff2a;
  rom[23262] = 16'hff2c;
  rom[23263] = 16'hf64b;
  rom[23264] = 16'hed49;
  rom[23265] = 16'hbb45;
  rom[23266] = 16'hbaa4;
  rom[23267] = 16'hd2e7;
  rom[23268] = 16'hca66;
  rom[23269] = 16'hcaa8;
  rom[23270] = 16'hb268;
  rom[23271] = 16'h7985;
  rom[23272] = 16'h92eb;
  rom[23273] = 16'he659;
  rom[23274] = 16'hffff;
  rom[23275] = 16'hffdf;
  rom[23276] = 16'hffff;
  rom[23277] = 16'hffff;
  rom[23278] = 16'hffbf;
  rom[23279] = 16'hffff;
  rom[23280] = 16'hffff;
  rom[23281] = 16'hffff;
  rom[23282] = 16'hffff;
  rom[23283] = 16'hffff;
  rom[23284] = 16'hffff;
  rom[23285] = 16'hffff;
  rom[23286] = 16'hffff;
  rom[23287] = 16'hffff;
  rom[23288] = 16'hffff;
  rom[23289] = 16'hffff;
  rom[23290] = 16'hffff;
  rom[23291] = 16'hffff;
  rom[23292] = 16'hffbd;
  rom[23293] = 16'hff7c;
  rom[23294] = 16'hff3a;
  rom[23295] = 16'hff1a;
  rom[23296] = 16'hfed9;
  rom[23297] = 16'hfefa;
  rom[23298] = 16'hfeda;
  rom[23299] = 16'hff3b;
  rom[23300] = 16'hff5c;
  rom[23301] = 16'hffbd;
  rom[23302] = 16'hffbe;
  rom[23303] = 16'hffff;
  rom[23304] = 16'hffff;
  rom[23305] = 16'hffff;
  rom[23306] = 16'hffff;
  rom[23307] = 16'hffff;
  rom[23308] = 16'hffff;
  rom[23309] = 16'hffff;
  rom[23310] = 16'hffff;
  rom[23311] = 16'hffff;
  rom[23312] = 16'hffff;
  rom[23313] = 16'hffff;
  rom[23314] = 16'hffde;
  rom[23315] = 16'hffdf;
  rom[23316] = 16'hffdf;
  rom[23317] = 16'hffdf;
  rom[23318] = 16'hf7bf;
  rom[23319] = 16'hffff;
  rom[23320] = 16'hf77c;
  rom[23321] = 16'hc4d2;
  rom[23322] = 16'h8a67;
  rom[23323] = 16'ha267;
  rom[23324] = 16'hc2c6;
  rom[23325] = 16'hcaa6;
  rom[23326] = 16'hcac5;
  rom[23327] = 16'hdb66;
  rom[23328] = 16'he426;
  rom[23329] = 16'hed08;
  rom[23330] = 16'hfe4a;
  rom[23331] = 16'hfecb;
  rom[23332] = 16'hfeeb;
  rom[23333] = 16'hfeeb;
  rom[23334] = 16'hff0b;
  rom[23335] = 16'hff2c;
  rom[23336] = 16'hef2d;
  rom[23337] = 16'hf70d;
  rom[23338] = 16'he68c;
  rom[23339] = 16'he62d;
  rom[23340] = 16'hc529;
  rom[23341] = 16'hb426;
  rom[23342] = 16'h9304;
  rom[23343] = 16'h7222;
  rom[23344] = 16'h69c1;
  rom[23345] = 16'h7203;
  rom[23346] = 16'h9ac8;
  rom[23347] = 16'hb34c;
  rom[23348] = 16'hbbad;
  rom[23349] = 16'hcc0e;
  rom[23350] = 16'hd42e;
  rom[23351] = 16'he4d2;
  rom[23352] = 16'he513;
  rom[23353] = 16'hed76;
  rom[23354] = 16'hed76;
  rom[23355] = 16'hf5f8;
  rom[23356] = 16'hf659;
  rom[23357] = 16'hfe99;
  rom[23358] = 16'hfeba;
  rom[23359] = 16'hfefb;
  rom[23360] = 16'hfeda;
  rom[23361] = 16'hff1c;
  rom[23362] = 16'hff3d;
  rom[23363] = 16'hff5d;
  rom[23364] = 16'hff3c;
  rom[23365] = 16'hff1c;
  rom[23366] = 16'hfedb;
  rom[23367] = 16'hfedb;
  rom[23368] = 16'hfedb;
  rom[23369] = 16'hfe7a;
  rom[23370] = 16'hfe18;
  rom[23371] = 16'hfdf7;
  rom[23372] = 16'hedb5;
  rom[23373] = 16'hed34;
  rom[23374] = 16'he471;
  rom[23375] = 16'hcc51;
  rom[23376] = 16'he678;
  rom[23377] = 16'hfffe;
  rom[23378] = 16'hffff;
  rom[23379] = 16'hffff;
  rom[23380] = 16'hffff;
  rom[23381] = 16'hffff;
  rom[23382] = 16'hffff;
  rom[23383] = 16'hffff;
  rom[23384] = 16'hffff;
  rom[23385] = 16'hffff;
  rom[23386] = 16'hffff;
  rom[23387] = 16'hffff;
  rom[23388] = 16'hffff;
  rom[23389] = 16'hffff;
  rom[23390] = 16'hffff;
  rom[23391] = 16'hffff;
  rom[23392] = 16'hffff;
  rom[23393] = 16'hffff;
  rom[23394] = 16'hffff;
  rom[23395] = 16'hffff;
  rom[23396] = 16'hffff;
  rom[23397] = 16'hffff;
  rom[23398] = 16'hffff;
  rom[23399] = 16'hffff;
  rom[23400] = 16'hffff;
  rom[23401] = 16'hffff;
  rom[23402] = 16'hffff;
  rom[23403] = 16'hffff;
  rom[23404] = 16'hffff;
  rom[23405] = 16'hffff;
  rom[23406] = 16'hffff;
  rom[23407] = 16'hffff;
  rom[23408] = 16'hffff;
  rom[23409] = 16'hffff;
  rom[23410] = 16'hffff;
  rom[23411] = 16'hffff;
  rom[23412] = 16'hffff;
  rom[23413] = 16'hffff;
  rom[23414] = 16'hffff;
  rom[23415] = 16'hffff;
  rom[23416] = 16'hffff;
  rom[23417] = 16'hffff;
  rom[23418] = 16'hffff;
  rom[23419] = 16'hffff;
  rom[23420] = 16'hffff;
  rom[23421] = 16'hffff;
  rom[23422] = 16'hffff;
  rom[23423] = 16'hffff;
  rom[23424] = 16'hffff;
  rom[23425] = 16'hffff;
  rom[23426] = 16'hffff;
  rom[23427] = 16'hffff;
  rom[23428] = 16'hffff;
  rom[23429] = 16'hffff;
  rom[23430] = 16'hffff;
  rom[23431] = 16'hffff;
  rom[23432] = 16'hffff;
  rom[23433] = 16'hffff;
  rom[23434] = 16'hffff;
  rom[23435] = 16'hffff;
  rom[23436] = 16'hffff;
  rom[23437] = 16'hffff;
  rom[23438] = 16'hffff;
  rom[23439] = 16'hffff;
  rom[23440] = 16'hffff;
  rom[23441] = 16'hffdf;
  rom[23442] = 16'hffdf;
  rom[23443] = 16'hffff;
  rom[23444] = 16'hffff;
  rom[23445] = 16'hffbf;
  rom[23446] = 16'hff9e;
  rom[23447] = 16'had11;
  rom[23448] = 16'h62a4;
  rom[23449] = 16'h83c5;
  rom[23450] = 16'he68d;
  rom[23451] = 16'hff2c;
  rom[23452] = 16'hff4b;
  rom[23453] = 16'hf6e9;
  rom[23454] = 16'hff2a;
  rom[23455] = 16'hfee9;
  rom[23456] = 16'hff08;
  rom[23457] = 16'hff09;
  rom[23458] = 16'hff2a;
  rom[23459] = 16'hff09;
  rom[23460] = 16'hff4b;
  rom[23461] = 16'hf70a;
  rom[23462] = 16'hfeea;
  rom[23463] = 16'hff0c;
  rom[23464] = 16'hfecc;
  rom[23465] = 16'hfdaa;
  rom[23466] = 16'hd3e5;
  rom[23467] = 16'hc303;
  rom[23468] = 16'hd2e6;
  rom[23469] = 16'hca87;
  rom[23470] = 16'hca67;
  rom[23471] = 16'hba48;
  rom[23472] = 16'h99a6;
  rom[23473] = 16'h9aaa;
  rom[23474] = 16'hd595;
  rom[23475] = 16'hff9d;
  rom[23476] = 16'hffff;
  rom[23477] = 16'hffff;
  rom[23478] = 16'hffff;
  rom[23479] = 16'hffff;
  rom[23480] = 16'hffff;
  rom[23481] = 16'hffff;
  rom[23482] = 16'hffff;
  rom[23483] = 16'hffff;
  rom[23484] = 16'hffff;
  rom[23485] = 16'hffff;
  rom[23486] = 16'hffff;
  rom[23487] = 16'hffff;
  rom[23488] = 16'hffff;
  rom[23489] = 16'hffff;
  rom[23490] = 16'hffff;
  rom[23491] = 16'hffff;
  rom[23492] = 16'hffff;
  rom[23493] = 16'hffbe;
  rom[23494] = 16'hffde;
  rom[23495] = 16'hfffe;
  rom[23496] = 16'hffff;
  rom[23497] = 16'hffff;
  rom[23498] = 16'hffff;
  rom[23499] = 16'hffff;
  rom[23500] = 16'hffff;
  rom[23501] = 16'hffff;
  rom[23502] = 16'hffff;
  rom[23503] = 16'hffff;
  rom[23504] = 16'hffff;
  rom[23505] = 16'hffff;
  rom[23506] = 16'hffff;
  rom[23507] = 16'hffff;
  rom[23508] = 16'hffff;
  rom[23509] = 16'hffff;
  rom[23510] = 16'hffff;
  rom[23511] = 16'hffff;
  rom[23512] = 16'hffff;
  rom[23513] = 16'hfffe;
  rom[23514] = 16'hffff;
  rom[23515] = 16'hffdf;
  rom[23516] = 16'hffff;
  rom[23517] = 16'hffdf;
  rom[23518] = 16'hffff;
  rom[23519] = 16'hf77c;
  rom[23520] = 16'ha42f;
  rom[23521] = 16'h7a25;
  rom[23522] = 16'haa87;
  rom[23523] = 16'hc2e7;
  rom[23524] = 16'hc2c4;
  rom[23525] = 16'hd387;
  rom[23526] = 16'hec48;
  rom[23527] = 16'hfd6a;
  rom[23528] = 16'hfe4a;
  rom[23529] = 16'hfeca;
  rom[23530] = 16'hff4b;
  rom[23531] = 16'hf74b;
  rom[23532] = 16'hf72c;
  rom[23533] = 16'hff0b;
  rom[23534] = 16'hff0b;
  rom[23535] = 16'hf6ea;
  rom[23536] = 16'hef2a;
  rom[23537] = 16'hef09;
  rom[23538] = 16'hff6c;
  rom[23539] = 16'hff4c;
  rom[23540] = 16'hff6e;
  rom[23541] = 16'hf70d;
  rom[23542] = 16'hfece;
  rom[23543] = 16'he5eb;
  rom[23544] = 16'hc487;
  rom[23545] = 16'h8ae2;
  rom[23546] = 16'h71c1;
  rom[23547] = 16'h7181;
  rom[23548] = 16'h89e4;
  rom[23549] = 16'ha266;
  rom[23550] = 16'hd32a;
  rom[23551] = 16'hc288;
  rom[23552] = 16'hc289;
  rom[23553] = 16'hca88;
  rom[23554] = 16'hcaca;
  rom[23555] = 16'hd30c;
  rom[23556] = 16'hdb4d;
  rom[23557] = 16'hd36d;
  rom[23558] = 16'he3ef;
  rom[23559] = 16'hdc0e;
  rom[23560] = 16'hdc0f;
  rom[23561] = 16'hdc2f;
  rom[23562] = 16'hec91;
  rom[23563] = 16'hec91;
  rom[23564] = 16'hec92;
  rom[23565] = 16'he450;
  rom[23566] = 16'he3ef;
  rom[23567] = 16'hdb8e;
  rom[23568] = 16'hebae;
  rom[23569] = 16'heb4d;
  rom[23570] = 16'he32d;
  rom[23571] = 16'hdb0b;
  rom[23572] = 16'hd2ca;
  rom[23573] = 16'hca68;
  rom[23574] = 16'hca29;
  rom[23575] = 16'hcb2c;
  rom[23576] = 16'hfe99;
  rom[23577] = 16'hfffe;
  rom[23578] = 16'hffff;
  rom[23579] = 16'hffff;
  rom[23580] = 16'hffff;
  rom[23581] = 16'hffff;
  rom[23582] = 16'hffff;
  rom[23583] = 16'hffff;
  rom[23584] = 16'hffff;
  rom[23585] = 16'hffff;
  rom[23586] = 16'hffff;
  rom[23587] = 16'hffff;
  rom[23588] = 16'hffff;
  rom[23589] = 16'hffff;
  rom[23590] = 16'hffff;
  rom[23591] = 16'hffff;
  rom[23592] = 16'hffff;
  rom[23593] = 16'hffff;
  rom[23594] = 16'hffff;
  rom[23595] = 16'hffff;
  rom[23596] = 16'hffff;
  rom[23597] = 16'hffff;
  rom[23598] = 16'hffff;
  rom[23599] = 16'hffff;
  rom[23600] = 16'hffff;
  rom[23601] = 16'hffff;
  rom[23602] = 16'hffff;
  rom[23603] = 16'hffff;
  rom[23604] = 16'hffff;
  rom[23605] = 16'hffff;
  rom[23606] = 16'hffff;
  rom[23607] = 16'hffff;
  rom[23608] = 16'hffff;
  rom[23609] = 16'hffff;
  rom[23610] = 16'hffff;
  rom[23611] = 16'hffff;
  rom[23612] = 16'hffdf;
  rom[23613] = 16'hffff;
  rom[23614] = 16'hffff;
  rom[23615] = 16'hffff;
  rom[23616] = 16'hffff;
  rom[23617] = 16'hffff;
  rom[23618] = 16'hffff;
  rom[23619] = 16'hffff;
  rom[23620] = 16'hffff;
  rom[23621] = 16'hffff;
  rom[23622] = 16'hffff;
  rom[23623] = 16'hffff;
  rom[23624] = 16'hffff;
  rom[23625] = 16'hffff;
  rom[23626] = 16'hffff;
  rom[23627] = 16'hffff;
  rom[23628] = 16'hffff;
  rom[23629] = 16'hffff;
  rom[23630] = 16'hffff;
  rom[23631] = 16'hffff;
  rom[23632] = 16'hffff;
  rom[23633] = 16'hffff;
  rom[23634] = 16'hfffe;
  rom[23635] = 16'hffff;
  rom[23636] = 16'hffdf;
  rom[23637] = 16'hffff;
  rom[23638] = 16'hffff;
  rom[23639] = 16'hffff;
  rom[23640] = 16'hffff;
  rom[23641] = 16'hffdf;
  rom[23642] = 16'hffdf;
  rom[23643] = 16'hffff;
  rom[23644] = 16'hffff;
  rom[23645] = 16'hffdf;
  rom[23646] = 16'hff9e;
  rom[23647] = 16'hff5c;
  rom[23648] = 16'hd593;
  rom[23649] = 16'h7a23;
  rom[23650] = 16'h7a61;
  rom[23651] = 16'hbc87;
  rom[23652] = 16'hf66c;
  rom[23653] = 16'hfecc;
  rom[23654] = 16'hf6e9;
  rom[23655] = 16'hff6a;
  rom[23656] = 16'hff28;
  rom[23657] = 16'hff09;
  rom[23658] = 16'hf709;
  rom[23659] = 16'hff0a;
  rom[23660] = 16'hff2a;
  rom[23661] = 16'hff2a;
  rom[23662] = 16'hf70a;
  rom[23663] = 16'hf72a;
  rom[23664] = 16'hff0a;
  rom[23665] = 16'hfeeb;
  rom[23666] = 16'hfe49;
  rom[23667] = 16'hfd89;
  rom[23668] = 16'he448;
  rom[23669] = 16'hd325;
  rom[23670] = 16'hc284;
  rom[23671] = 16'hd2a7;
  rom[23672] = 16'hc287;
  rom[23673] = 16'haa68;
  rom[23674] = 16'h8a67;
  rom[23675] = 16'hb470;
  rom[23676] = 16'hf71b;
  rom[23677] = 16'hffde;
  rom[23678] = 16'hffff;
  rom[23679] = 16'hffff;
  rom[23680] = 16'hffff;
  rom[23681] = 16'hffff;
  rom[23682] = 16'hffff;
  rom[23683] = 16'hffff;
  rom[23684] = 16'hffff;
  rom[23685] = 16'hffff;
  rom[23686] = 16'hffff;
  rom[23687] = 16'hffff;
  rom[23688] = 16'hffff;
  rom[23689] = 16'hffff;
  rom[23690] = 16'hffff;
  rom[23691] = 16'hffff;
  rom[23692] = 16'hffdf;
  rom[23693] = 16'hffff;
  rom[23694] = 16'hffff;
  rom[23695] = 16'hffff;
  rom[23696] = 16'hffff;
  rom[23697] = 16'hffff;
  rom[23698] = 16'hffff;
  rom[23699] = 16'hffff;
  rom[23700] = 16'hffff;
  rom[23701] = 16'hffff;
  rom[23702] = 16'hffdf;
  rom[23703] = 16'hffff;
  rom[23704] = 16'hffff;
  rom[23705] = 16'hffff;
  rom[23706] = 16'hffff;
  rom[23707] = 16'hffff;
  rom[23708] = 16'hffff;
  rom[23709] = 16'hffff;
  rom[23710] = 16'hfffe;
  rom[23711] = 16'hffff;
  rom[23712] = 16'hfffe;
  rom[23713] = 16'hffff;
  rom[23714] = 16'hffff;
  rom[23715] = 16'hffff;
  rom[23716] = 16'hffff;
  rom[23717] = 16'hffbe;
  rom[23718] = 16'hcdd6;
  rom[23719] = 16'h830a;
  rom[23720] = 16'h82a6;
  rom[23721] = 16'ha2e6;
  rom[23722] = 16'hc345;
  rom[23723] = 16'hdbc6;
  rom[23724] = 16'hf509;
  rom[23725] = 16'hfdec;
  rom[23726] = 16'hfe4c;
  rom[23727] = 16'hfeab;
  rom[23728] = 16'hfeea;
  rom[23729] = 16'hff08;
  rom[23730] = 16'hf728;
  rom[23731] = 16'hf74a;
  rom[23732] = 16'hf70b;
  rom[23733] = 16'hf70b;
  rom[23734] = 16'hf6c9;
  rom[23735] = 16'hff2a;
  rom[23736] = 16'hf729;
  rom[23737] = 16'hff4a;
  rom[23738] = 16'hef4a;
  rom[23739] = 16'hef29;
  rom[23740] = 16'hef09;
  rom[23741] = 16'hf72b;
  rom[23742] = 16'hf6ea;
  rom[23743] = 16'hff0b;
  rom[23744] = 16'hfeab;
  rom[23745] = 16'hfe8c;
  rom[23746] = 16'hddca;
  rom[23747] = 16'hbc66;
  rom[23748] = 16'h8aa2;
  rom[23749] = 16'h79a1;
  rom[23750] = 16'h8982;
  rom[23751] = 16'hb246;
  rom[23752] = 16'hc267;
  rom[23753] = 16'hd2a8;
  rom[23754] = 16'hd266;
  rom[23755] = 16'he288;
  rom[23756] = 16'hda27;
  rom[23757] = 16'hda27;
  rom[23758] = 16'hda47;
  rom[23759] = 16'he268;
  rom[23760] = 16'hda48;
  rom[23761] = 16'hda68;
  rom[23762] = 16'hd268;
  rom[23763] = 16'hd268;
  rom[23764] = 16'hca47;
  rom[23765] = 16'hd248;
  rom[23766] = 16'hda48;
  rom[23767] = 16'he248;
  rom[23768] = 16'he228;
  rom[23769] = 16'hf249;
  rom[23770] = 16'he228;
  rom[23771] = 16'he227;
  rom[23772] = 16'hda06;
  rom[23773] = 16'hea28;
  rom[23774] = 16'hda07;
  rom[23775] = 16'hdacb;
  rom[23776] = 16'hfe78;
  rom[23777] = 16'hffdd;
  rom[23778] = 16'hffde;
  rom[23779] = 16'hffff;
  rom[23780] = 16'hffff;
  rom[23781] = 16'hffff;
  rom[23782] = 16'hffff;
  rom[23783] = 16'hffff;
  rom[23784] = 16'hffff;
  rom[23785] = 16'hffff;
  rom[23786] = 16'hffff;
  rom[23787] = 16'hffff;
  rom[23788] = 16'hffff;
  rom[23789] = 16'hffff;
  rom[23790] = 16'hffff;
  rom[23791] = 16'hffff;
  rom[23792] = 16'hffff;
  rom[23793] = 16'hffff;
  rom[23794] = 16'hffff;
  rom[23795] = 16'hffff;
  rom[23796] = 16'hffff;
  rom[23797] = 16'hffff;
  rom[23798] = 16'hffff;
  rom[23799] = 16'hffff;
  rom[23800] = 16'hffff;
  rom[23801] = 16'hffff;
  rom[23802] = 16'hffff;
  rom[23803] = 16'hffff;
  rom[23804] = 16'hffff;
  rom[23805] = 16'hffff;
  rom[23806] = 16'hffff;
  rom[23807] = 16'hffff;
  rom[23808] = 16'hffff;
  rom[23809] = 16'hffff;
  rom[23810] = 16'hffff;
  rom[23811] = 16'hffff;
  rom[23812] = 16'hffff;
  rom[23813] = 16'hffff;
  rom[23814] = 16'hffff;
  rom[23815] = 16'hffff;
  rom[23816] = 16'hffff;
  rom[23817] = 16'hffff;
  rom[23818] = 16'hffff;
  rom[23819] = 16'hffff;
  rom[23820] = 16'hffff;
  rom[23821] = 16'hffff;
  rom[23822] = 16'hffff;
  rom[23823] = 16'hffff;
  rom[23824] = 16'hffff;
  rom[23825] = 16'hffff;
  rom[23826] = 16'hffff;
  rom[23827] = 16'hffff;
  rom[23828] = 16'hffff;
  rom[23829] = 16'hffff;
  rom[23830] = 16'hffff;
  rom[23831] = 16'hffff;
  rom[23832] = 16'hffff;
  rom[23833] = 16'hffff;
  rom[23834] = 16'hfffe;
  rom[23835] = 16'hfffe;
  rom[23836] = 16'hffff;
  rom[23837] = 16'hffff;
  rom[23838] = 16'hffff;
  rom[23839] = 16'hffff;
  rom[23840] = 16'hffff;
  rom[23841] = 16'hffff;
  rom[23842] = 16'hffff;
  rom[23843] = 16'hffff;
  rom[23844] = 16'hffff;
  rom[23845] = 16'hffff;
  rom[23846] = 16'hff9e;
  rom[23847] = 16'hf5f7;
  rom[23848] = 16'hbb4b;
  rom[23849] = 16'hc32a;
  rom[23850] = 16'haa25;
  rom[23851] = 16'h6900;
  rom[23852] = 16'ha346;
  rom[23853] = 16'hd56a;
  rom[23854] = 16'hff4e;
  rom[23855] = 16'he6a8;
  rom[23856] = 16'hf709;
  rom[23857] = 16'hf749;
  rom[23858] = 16'hff29;
  rom[23859] = 16'hff6b;
  rom[23860] = 16'hf709;
  rom[23861] = 16'hf709;
  rom[23862] = 16'hff6a;
  rom[23863] = 16'hf708;
  rom[23864] = 16'hff6b;
  rom[23865] = 16'hff08;
  rom[23866] = 16'hfee9;
  rom[23867] = 16'hff0b;
  rom[23868] = 16'hfeac;
  rom[23869] = 16'hfdca;
  rom[23870] = 16'hec88;
  rom[23871] = 16'hdba6;
  rom[23872] = 16'hd2e5;
  rom[23873] = 16'hba65;
  rom[23874] = 16'hc349;
  rom[23875] = 16'h79c4;
  rom[23876] = 16'h7a88;
  rom[23877] = 16'hde57;
  rom[23878] = 16'hffde;
  rom[23879] = 16'hffbd;
  rom[23880] = 16'hffff;
  rom[23881] = 16'hffff;
  rom[23882] = 16'hffff;
  rom[23883] = 16'hffff;
  rom[23884] = 16'hffff;
  rom[23885] = 16'hffff;
  rom[23886] = 16'hfffe;
  rom[23887] = 16'hffff;
  rom[23888] = 16'hffff;
  rom[23889] = 16'hffff;
  rom[23890] = 16'hffff;
  rom[23891] = 16'hffff;
  rom[23892] = 16'hffff;
  rom[23893] = 16'hffff;
  rom[23894] = 16'hffff;
  rom[23895] = 16'hffff;
  rom[23896] = 16'hffff;
  rom[23897] = 16'hffff;
  rom[23898] = 16'hffff;
  rom[23899] = 16'hffff;
  rom[23900] = 16'hffff;
  rom[23901] = 16'hffff;
  rom[23902] = 16'hffde;
  rom[23903] = 16'hffff;
  rom[23904] = 16'hffff;
  rom[23905] = 16'hffff;
  rom[23906] = 16'hffff;
  rom[23907] = 16'hffff;
  rom[23908] = 16'hffff;
  rom[23909] = 16'hffff;
  rom[23910] = 16'hffff;
  rom[23911] = 16'hffde;
  rom[23912] = 16'hffff;
  rom[23913] = 16'hffff;
  rom[23914] = 16'hfffe;
  rom[23915] = 16'hfffe;
  rom[23916] = 16'hff7c;
  rom[23917] = 16'hbcd0;
  rom[23918] = 16'h7224;
  rom[23919] = 16'h92e6;
  rom[23920] = 16'hab46;
  rom[23921] = 16'hc3e6;
  rom[23922] = 16'hf589;
  rom[23923] = 16'hfe6b;
  rom[23924] = 16'hfeac;
  rom[23925] = 16'hfe6a;
  rom[23926] = 16'hfecb;
  rom[23927] = 16'hff0a;
  rom[23928] = 16'hff0a;
  rom[23929] = 16'hff48;
  rom[23930] = 16'hff69;
  rom[23931] = 16'hff29;
  rom[23932] = 16'hff4b;
  rom[23933] = 16'hff2a;
  rom[23934] = 16'hff4a;
  rom[23935] = 16'hff28;
  rom[23936] = 16'hff29;
  rom[23937] = 16'heee7;
  rom[23938] = 16'hff69;
  rom[23939] = 16'hff8a;
  rom[23940] = 16'hff69;
  rom[23941] = 16'hf748;
  rom[23942] = 16'hff6a;
  rom[23943] = 16'hff6a;
  rom[23944] = 16'hff2b;
  rom[23945] = 16'hf70a;
  rom[23946] = 16'hf70b;
  rom[23947] = 16'heeaa;
  rom[23948] = 16'hff2e;
  rom[23949] = 16'hdd6b;
  rom[23950] = 16'ha324;
  rom[23951] = 16'h6920;
  rom[23952] = 16'h8941;
  rom[23953] = 16'hb246;
  rom[23954] = 16'hd2a7;
  rom[23955] = 16'hda67;
  rom[23956] = 16'hea68;
  rom[23957] = 16'hea26;
  rom[23958] = 16'hf207;
  rom[23959] = 16'hea07;
  rom[23960] = 16'hf207;
  rom[23961] = 16'he1e6;
  rom[23962] = 16'hf289;
  rom[23963] = 16'hea68;
  rom[23964] = 16'he268;
  rom[23965] = 16'he247;
  rom[23966] = 16'hea47;
  rom[23967] = 16'hea06;
  rom[23968] = 16'he9c6;
  rom[23969] = 16'hf1c6;
  rom[23970] = 16'hf227;
  rom[23971] = 16'hf246;
  rom[23972] = 16'hf226;
  rom[23973] = 16'hf206;
  rom[23974] = 16'he9e7;
  rom[23975] = 16'he2eb;
  rom[23976] = 16'hfe99;
  rom[23977] = 16'hfffe;
  rom[23978] = 16'hffff;
  rom[23979] = 16'hffff;
  rom[23980] = 16'hffff;
  rom[23981] = 16'hffff;
  rom[23982] = 16'hffff;
  rom[23983] = 16'hffff;
  rom[23984] = 16'hffff;
  rom[23985] = 16'hffff;
  rom[23986] = 16'hffff;
  rom[23987] = 16'hffff;
  rom[23988] = 16'hffff;
  rom[23989] = 16'hffff;
  rom[23990] = 16'hffff;
  rom[23991] = 16'hffff;
  rom[23992] = 16'hffff;
  rom[23993] = 16'hffff;
  rom[23994] = 16'hffff;
  rom[23995] = 16'hffff;
  rom[23996] = 16'hffff;
  rom[23997] = 16'hffff;
  rom[23998] = 16'hffff;
  rom[23999] = 16'hffff;
  rom[24000] = 16'hffff;
  rom[24001] = 16'hffff;
  rom[24002] = 16'hffff;
  rom[24003] = 16'hffff;
  rom[24004] = 16'hffdf;
  rom[24005] = 16'hffff;
  rom[24006] = 16'hffdf;
  rom[24007] = 16'hffff;
  rom[24008] = 16'hffff;
  rom[24009] = 16'hffff;
  rom[24010] = 16'hff7d;
  rom[24011] = 16'hffbf;
  rom[24012] = 16'hffdf;
  rom[24013] = 16'hffff;
  rom[24014] = 16'hffff;
  rom[24015] = 16'hffff;
  rom[24016] = 16'hffff;
  rom[24017] = 16'hffff;
  rom[24018] = 16'hffff;
  rom[24019] = 16'hffff;
  rom[24020] = 16'hffff;
  rom[24021] = 16'hffff;
  rom[24022] = 16'hffff;
  rom[24023] = 16'hffff;
  rom[24024] = 16'hffff;
  rom[24025] = 16'hffff;
  rom[24026] = 16'hffff;
  rom[24027] = 16'hffff;
  rom[24028] = 16'hffff;
  rom[24029] = 16'hffff;
  rom[24030] = 16'hffff;
  rom[24031] = 16'hffff;
  rom[24032] = 16'hffff;
  rom[24033] = 16'hffff;
  rom[24034] = 16'hffff;
  rom[24035] = 16'hffff;
  rom[24036] = 16'hffdf;
  rom[24037] = 16'hffff;
  rom[24038] = 16'hffff;
  rom[24039] = 16'hffff;
  rom[24040] = 16'hffff;
  rom[24041] = 16'hffff;
  rom[24042] = 16'hffff;
  rom[24043] = 16'hffde;
  rom[24044] = 16'hffdd;
  rom[24045] = 16'hff5b;
  rom[24046] = 16'hed94;
  rom[24047] = 16'hd38d;
  rom[24048] = 16'hd288;
  rom[24049] = 16'hd248;
  rom[24050] = 16'hd248;
  rom[24051] = 16'hba47;
  rom[24052] = 16'h7962;
  rom[24053] = 16'h79e1;
  rom[24054] = 16'ha405;
  rom[24055] = 16'he68d;
  rom[24056] = 16'hf72c;
  rom[24057] = 16'hf70b;
  rom[24058] = 16'hf729;
  rom[24059] = 16'hf729;
  rom[24060] = 16'hf728;
  rom[24061] = 16'hff48;
  rom[24062] = 16'hf728;
  rom[24063] = 16'hff49;
  rom[24064] = 16'hf729;
  rom[24065] = 16'hff29;
  rom[24066] = 16'hf709;
  rom[24067] = 16'hff09;
  rom[24068] = 16'hfee9;
  rom[24069] = 16'hfeca;
  rom[24070] = 16'hfeaa;
  rom[24071] = 16'hfde9;
  rom[24072] = 16'he4e7;
  rom[24073] = 16'hdc27;
  rom[24074] = 16'hcb46;
  rom[24075] = 16'hbb08;
  rom[24076] = 16'h8a65;
  rom[24077] = 16'h7a67;
  rom[24078] = 16'h940d;
  rom[24079] = 16'hce17;
  rom[24080] = 16'hf77c;
  rom[24081] = 16'hffff;
  rom[24082] = 16'hffff;
  rom[24083] = 16'hffff;
  rom[24084] = 16'hffdf;
  rom[24085] = 16'hffff;
  rom[24086] = 16'hfffe;
  rom[24087] = 16'hffff;
  rom[24088] = 16'hfffe;
  rom[24089] = 16'hffff;
  rom[24090] = 16'hffff;
  rom[24091] = 16'hffff;
  rom[24092] = 16'hffff;
  rom[24093] = 16'hffff;
  rom[24094] = 16'hffff;
  rom[24095] = 16'hffff;
  rom[24096] = 16'hffff;
  rom[24097] = 16'hffff;
  rom[24098] = 16'hffff;
  rom[24099] = 16'hffff;
  rom[24100] = 16'hffff;
  rom[24101] = 16'hffff;
  rom[24102] = 16'hffff;
  rom[24103] = 16'hffff;
  rom[24104] = 16'hfffe;
  rom[24105] = 16'hffff;
  rom[24106] = 16'hffff;
  rom[24107] = 16'hffff;
  rom[24108] = 16'hf7ff;
  rom[24109] = 16'hffff;
  rom[24110] = 16'hffdf;
  rom[24111] = 16'hffff;
  rom[24112] = 16'hfffe;
  rom[24113] = 16'hfffe;
  rom[24114] = 16'he6f9;
  rom[24115] = 16'hb511;
  rom[24116] = 16'h6aa5;
  rom[24117] = 16'h7a84;
  rom[24118] = 16'hb3a7;
  rom[24119] = 16'hcc69;
  rom[24120] = 16'hedab;
  rom[24121] = 16'hfe6b;
  rom[24122] = 16'hfec9;
  rom[24123] = 16'hff29;
  rom[24124] = 16'hff28;
  rom[24125] = 16'hff2a;
  rom[24126] = 16'hff2a;
  rom[24127] = 16'hff2b;
  rom[24128] = 16'hf6e9;
  rom[24129] = 16'hff29;
  rom[24130] = 16'hfee8;
  rom[24131] = 16'hff09;
  rom[24132] = 16'hf708;
  rom[24133] = 16'hff28;
  rom[24134] = 16'hff49;
  rom[24135] = 16'hf707;
  rom[24136] = 16'hff48;
  rom[24137] = 16'hff49;
  rom[24138] = 16'hf708;
  rom[24139] = 16'hff08;
  rom[24140] = 16'hff08;
  rom[24141] = 16'hf708;
  rom[24142] = 16'hff29;
  rom[24143] = 16'hf709;
  rom[24144] = 16'hef09;
  rom[24145] = 16'hf74a;
  rom[24146] = 16'hf70a;
  rom[24147] = 16'hff4b;
  rom[24148] = 16'hf6ea;
  rom[24149] = 16'hfeec;
  rom[24150] = 16'hf6ac;
  rom[24151] = 16'hd58b;
  rom[24152] = 16'h9b65;
  rom[24153] = 16'h71e2;
  rom[24154] = 16'h89a3;
  rom[24155] = 16'hb266;
  rom[24156] = 16'hca66;
  rom[24157] = 16'hda67;
  rom[24158] = 16'hea07;
  rom[24159] = 16'hf1e7;
  rom[24160] = 16'hf207;
  rom[24161] = 16'hf227;
  rom[24162] = 16'hea06;
  rom[24163] = 16'hea47;
  rom[24164] = 16'he226;
  rom[24165] = 16'he247;
  rom[24166] = 16'he247;
  rom[24167] = 16'hea46;
  rom[24168] = 16'he226;
  rom[24169] = 16'hf226;
  rom[24170] = 16'he206;
  rom[24171] = 16'he245;
  rom[24172] = 16'he225;
  rom[24173] = 16'hf246;
  rom[24174] = 16'he206;
  rom[24175] = 16'he30b;
  rom[24176] = 16'hfed9;
  rom[24177] = 16'hfffe;
  rom[24178] = 16'hffff;
  rom[24179] = 16'hffff;
  rom[24180] = 16'hffff;
  rom[24181] = 16'hffff;
  rom[24182] = 16'hffff;
  rom[24183] = 16'hffff;
  rom[24184] = 16'hffff;
  rom[24185] = 16'hffff;
  rom[24186] = 16'hffff;
  rom[24187] = 16'hffff;
  rom[24188] = 16'hffff;
  rom[24189] = 16'hffff;
  rom[24190] = 16'hffff;
  rom[24191] = 16'hffff;
  rom[24192] = 16'hffff;
  rom[24193] = 16'hffff;
  rom[24194] = 16'hffff;
  rom[24195] = 16'hffff;
  rom[24196] = 16'hffff;
  rom[24197] = 16'hffff;
  rom[24198] = 16'hffff;
  rom[24199] = 16'hffff;
  rom[24200] = 16'hffff;
  rom[24201] = 16'hffff;
  rom[24202] = 16'hffff;
  rom[24203] = 16'hffff;
  rom[24204] = 16'hffff;
  rom[24205] = 16'hffff;
  rom[24206] = 16'hffff;
  rom[24207] = 16'hffff;
  rom[24208] = 16'hffff;
  rom[24209] = 16'hfffe;
  rom[24210] = 16'hdd75;
  rom[24211] = 16'hf67a;
  rom[24212] = 16'hff7e;
  rom[24213] = 16'hffde;
  rom[24214] = 16'hffff;
  rom[24215] = 16'hffff;
  rom[24216] = 16'hffff;
  rom[24217] = 16'hffff;
  rom[24218] = 16'hffff;
  rom[24219] = 16'hffff;
  rom[24220] = 16'hffff;
  rom[24221] = 16'hffff;
  rom[24222] = 16'hffff;
  rom[24223] = 16'hffff;
  rom[24224] = 16'hffff;
  rom[24225] = 16'hffff;
  rom[24226] = 16'hffff;
  rom[24227] = 16'hffff;
  rom[24228] = 16'hffff;
  rom[24229] = 16'hffff;
  rom[24230] = 16'hffff;
  rom[24231] = 16'hffff;
  rom[24232] = 16'hffff;
  rom[24233] = 16'hffff;
  rom[24234] = 16'hffff;
  rom[24235] = 16'hffff;
  rom[24236] = 16'hffff;
  rom[24237] = 16'hffff;
  rom[24238] = 16'hffff;
  rom[24239] = 16'hffff;
  rom[24240] = 16'hffff;
  rom[24241] = 16'hffff;
  rom[24242] = 16'hffbe;
  rom[24243] = 16'hff7d;
  rom[24244] = 16'hfef9;
  rom[24245] = 16'hdc8f;
  rom[24246] = 16'hcb2a;
  rom[24247] = 16'hda88;
  rom[24248] = 16'hea48;
  rom[24249] = 16'hea27;
  rom[24250] = 16'he228;
  rom[24251] = 16'hd248;
  rom[24252] = 16'hc267;
  rom[24253] = 16'ha245;
  rom[24254] = 16'h7161;
  rom[24255] = 16'h7202;
  rom[24256] = 16'hc4a8;
  rom[24257] = 16'hfeee;
  rom[24258] = 16'hf6cc;
  rom[24259] = 16'hff6c;
  rom[24260] = 16'hf709;
  rom[24261] = 16'hef07;
  rom[24262] = 16'hff6a;
  rom[24263] = 16'hf6c8;
  rom[24264] = 16'hff0a;
  rom[24265] = 16'hff2a;
  rom[24266] = 16'hff2a;
  rom[24267] = 16'hf6e8;
  rom[24268] = 16'hff09;
  rom[24269] = 16'hff08;
  rom[24270] = 16'hff09;
  rom[24271] = 16'hff2a;
  rom[24272] = 16'hfeec;
  rom[24273] = 16'hfe4c;
  rom[24274] = 16'hfdac;
  rom[24275] = 16'hecca;
  rom[24276] = 16'hc429;
  rom[24277] = 16'h9b46;
  rom[24278] = 16'h8b46;
  rom[24279] = 16'h6aa6;
  rom[24280] = 16'h7329;
  rom[24281] = 16'hb552;
  rom[24282] = 16'hfffe;
  rom[24283] = 16'hffbe;
  rom[24284] = 16'hffff;
  rom[24285] = 16'hfffe;
  rom[24286] = 16'hffff;
  rom[24287] = 16'hffff;
  rom[24288] = 16'hffff;
  rom[24289] = 16'hffff;
  rom[24290] = 16'hffff;
  rom[24291] = 16'hffff;
  rom[24292] = 16'hffff;
  rom[24293] = 16'hffff;
  rom[24294] = 16'hffff;
  rom[24295] = 16'hffff;
  rom[24296] = 16'hffdf;
  rom[24297] = 16'hffff;
  rom[24298] = 16'hffff;
  rom[24299] = 16'hffff;
  rom[24300] = 16'hffff;
  rom[24301] = 16'hffff;
  rom[24302] = 16'hffff;
  rom[24303] = 16'hffdf;
  rom[24304] = 16'hffff;
  rom[24305] = 16'hffdf;
  rom[24306] = 16'hffff;
  rom[24307] = 16'hffff;
  rom[24308] = 16'hf7df;
  rom[24309] = 16'hffff;
  rom[24310] = 16'hffff;
  rom[24311] = 16'hfffe;
  rom[24312] = 16'hef19;
  rom[24313] = 16'h946d;
  rom[24314] = 16'h62a4;
  rom[24315] = 16'h8345;
  rom[24316] = 16'hbcc9;
  rom[24317] = 16'hdd6a;
  rom[24318] = 16'hfe2d;
  rom[24319] = 16'hfe8d;
  rom[24320] = 16'hfecc;
  rom[24321] = 16'hfeea;
  rom[24322] = 16'hff29;
  rom[24323] = 16'hf748;
  rom[24324] = 16'hff69;
  rom[24325] = 16'hff49;
  rom[24326] = 16'hff6a;
  rom[24327] = 16'heeea;
  rom[24328] = 16'hf70b;
  rom[24329] = 16'hf72c;
  rom[24330] = 16'hff0c;
  rom[24331] = 16'hff2c;
  rom[24332] = 16'hf6e9;
  rom[24333] = 16'hff4a;
  rom[24334] = 16'heee8;
  rom[24335] = 16'hff49;
  rom[24336] = 16'hf708;
  rom[24337] = 16'hf708;
  rom[24338] = 16'hff09;
  rom[24339] = 16'hff29;
  rom[24340] = 16'hff09;
  rom[24341] = 16'hff09;
  rom[24342] = 16'hff29;
  rom[24343] = 16'hff09;
  rom[24344] = 16'hff4a;
  rom[24345] = 16'hf729;
  rom[24346] = 16'hff2a;
  rom[24347] = 16'hff29;
  rom[24348] = 16'hff2a;
  rom[24349] = 16'hf729;
  rom[24350] = 16'hf72a;
  rom[24351] = 16'hf72c;
  rom[24352] = 16'hee8d;
  rom[24353] = 16'hcd6b;
  rom[24354] = 16'h9b25;
  rom[24355] = 16'h68e0;
  rom[24356] = 16'h99a3;
  rom[24357] = 16'hca87;
  rom[24358] = 16'he288;
  rom[24359] = 16'hda06;
  rom[24360] = 16'hea27;
  rom[24361] = 16'hea07;
  rom[24362] = 16'he9c7;
  rom[24363] = 16'hf227;
  rom[24364] = 16'hf247;
  rom[24365] = 16'he247;
  rom[24366] = 16'hea47;
  rom[24367] = 16'he226;
  rom[24368] = 16'hea46;
  rom[24369] = 16'hea26;
  rom[24370] = 16'hea47;
  rom[24371] = 16'hea46;
  rom[24372] = 16'hf246;
  rom[24373] = 16'he246;
  rom[24374] = 16'he288;
  rom[24375] = 16'hdb2c;
  rom[24376] = 16'hff5b;
  rom[24377] = 16'hffff;
  rom[24378] = 16'hffff;
  rom[24379] = 16'hffff;
  rom[24380] = 16'hffff;
  rom[24381] = 16'hffff;
  rom[24382] = 16'hffff;
  rom[24383] = 16'hffff;
  rom[24384] = 16'hffff;
  rom[24385] = 16'hffff;
  rom[24386] = 16'hffff;
  rom[24387] = 16'hffff;
  rom[24388] = 16'hffff;
  rom[24389] = 16'hffff;
  rom[24390] = 16'hffff;
  rom[24391] = 16'hffff;
  rom[24392] = 16'hffff;
  rom[24393] = 16'hffff;
  rom[24394] = 16'hffff;
  rom[24395] = 16'hffff;
  rom[24396] = 16'hffff;
  rom[24397] = 16'hffff;
  rom[24398] = 16'hffff;
  rom[24399] = 16'hffff;
  rom[24400] = 16'hffdf;
  rom[24401] = 16'hffff;
  rom[24402] = 16'hf7fe;
  rom[24403] = 16'hffff;
  rom[24404] = 16'hffff;
  rom[24405] = 16'hffff;
  rom[24406] = 16'hffdf;
  rom[24407] = 16'hffff;
  rom[24408] = 16'hf7ff;
  rom[24409] = 16'hfffe;
  rom[24410] = 16'hab6c;
  rom[24411] = 16'hcc0f;
  rom[24412] = 16'hfe17;
  rom[24413] = 16'hffbd;
  rom[24414] = 16'hffbd;
  rom[24415] = 16'hffff;
  rom[24416] = 16'hffff;
  rom[24417] = 16'hffff;
  rom[24418] = 16'hffff;
  rom[24419] = 16'hffff;
  rom[24420] = 16'hffff;
  rom[24421] = 16'hffff;
  rom[24422] = 16'hffff;
  rom[24423] = 16'hffff;
  rom[24424] = 16'hffff;
  rom[24425] = 16'hffff;
  rom[24426] = 16'hffff;
  rom[24427] = 16'hffff;
  rom[24428] = 16'hffff;
  rom[24429] = 16'hffff;
  rom[24430] = 16'hffff;
  rom[24431] = 16'hffff;
  rom[24432] = 16'hffff;
  rom[24433] = 16'hffff;
  rom[24434] = 16'hffff;
  rom[24435] = 16'hffff;
  rom[24436] = 16'hffdf;
  rom[24437] = 16'hffff;
  rom[24438] = 16'hfffe;
  rom[24439] = 16'hfffe;
  rom[24440] = 16'hffde;
  rom[24441] = 16'hff7d;
  rom[24442] = 16'hfeb9;
  rom[24443] = 16'hf554;
  rom[24444] = 16'hcb8c;
  rom[24445] = 16'hcac8;
  rom[24446] = 16'hd266;
  rom[24447] = 16'hea47;
  rom[24448] = 16'hf226;
  rom[24449] = 16'hf206;
  rom[24450] = 16'he225;
  rom[24451] = 16'hda47;
  rom[24452] = 16'he2a9;
  rom[24453] = 16'hca47;
  rom[24454] = 16'hc2a7;
  rom[24455] = 16'h99a3;
  rom[24456] = 16'h7141;
  rom[24457] = 16'h8a42;
  rom[24458] = 16'hdd6b;
  rom[24459] = 16'hf64c;
  rom[24460] = 16'hff2d;
  rom[24461] = 16'hff0b;
  rom[24462] = 16'hf6c9;
  rom[24463] = 16'hff4a;
  rom[24464] = 16'hff0a;
  rom[24465] = 16'hff2a;
  rom[24466] = 16'hf72a;
  rom[24467] = 16'hff2a;
  rom[24468] = 16'hff29;
  rom[24469] = 16'hff49;
  rom[24470] = 16'hf728;
  rom[24471] = 16'hf708;
  rom[24472] = 16'hff0a;
  rom[24473] = 16'hff2b;
  rom[24474] = 16'hfeab;
  rom[24475] = 16'hfe8c;
  rom[24476] = 16'hfeae;
  rom[24477] = 16'hfe4d;
  rom[24478] = 16'hddab;
  rom[24479] = 16'hbce9;
  rom[24480] = 16'h9408;
  rom[24481] = 16'h6aa4;
  rom[24482] = 16'h5285;
  rom[24483] = 16'h9ccf;
  rom[24484] = 16'hd656;
  rom[24485] = 16'hef3a;
  rom[24486] = 16'hffbc;
  rom[24487] = 16'hfffe;
  rom[24488] = 16'hffbe;
  rom[24489] = 16'hffff;
  rom[24490] = 16'hffdf;
  rom[24491] = 16'hffff;
  rom[24492] = 16'hffdf;
  rom[24493] = 16'hffff;
  rom[24494] = 16'hffff;
  rom[24495] = 16'hffff;
  rom[24496] = 16'hffdf;
  rom[24497] = 16'hffff;
  rom[24498] = 16'hffdf;
  rom[24499] = 16'hffff;
  rom[24500] = 16'hffff;
  rom[24501] = 16'hffff;
  rom[24502] = 16'hffff;
  rom[24503] = 16'hffdf;
  rom[24504] = 16'hffdf;
  rom[24505] = 16'hffbe;
  rom[24506] = 16'hffdf;
  rom[24507] = 16'hfffe;
  rom[24508] = 16'hf79c;
  rom[24509] = 16'he719;
  rom[24510] = 16'hc614;
  rom[24511] = 16'h942b;
  rom[24512] = 16'h62a3;
  rom[24513] = 16'h9407;
  rom[24514] = 16'hb52a;
  rom[24515] = 16'he66d;
  rom[24516] = 16'hf6cc;
  rom[24517] = 16'hfeec;
  rom[24518] = 16'hfeea;
  rom[24519] = 16'hfeea;
  rom[24520] = 16'hff0a;
  rom[24521] = 16'hff2a;
  rom[24522] = 16'hf729;
  rom[24523] = 16'hf729;
  rom[24524] = 16'heec7;
  rom[24525] = 16'hf6e8;
  rom[24526] = 16'hf728;
  rom[24527] = 16'hff6b;
  rom[24528] = 16'heecc;
  rom[24529] = 16'h8ba2;
  rom[24530] = 16'h93c4;
  rom[24531] = 16'he68e;
  rom[24532] = 16'heeec;
  rom[24533] = 16'hff4c;
  rom[24534] = 16'hf74a;
  rom[24535] = 16'hf729;
  rom[24536] = 16'hff49;
  rom[24537] = 16'hff29;
  rom[24538] = 16'hf709;
  rom[24539] = 16'hfee9;
  rom[24540] = 16'hfee9;
  rom[24541] = 16'hff29;
  rom[24542] = 16'hf6e8;
  rom[24543] = 16'hff29;
  rom[24544] = 16'hf729;
  rom[24545] = 16'hf729;
  rom[24546] = 16'hf709;
  rom[24547] = 16'hf729;
  rom[24548] = 16'hff29;
  rom[24549] = 16'hff09;
  rom[24550] = 16'hf6e8;
  rom[24551] = 16'hff4a;
  rom[24552] = 16'hf74c;
  rom[24553] = 16'hff2d;
  rom[24554] = 16'hf6ae;
  rom[24555] = 16'hccaa;
  rom[24556] = 16'h79e1;
  rom[24557] = 16'h8162;
  rom[24558] = 16'haa65;
  rom[24559] = 16'hcaa8;
  rom[24560] = 16'hd227;
  rom[24561] = 16'hea07;
  rom[24562] = 16'hfa28;
  rom[24563] = 16'hf1c6;
  rom[24564] = 16'hf1e6;
  rom[24565] = 16'hf206;
  rom[24566] = 16'hea26;
  rom[24567] = 16'hea46;
  rom[24568] = 16'hea46;
  rom[24569] = 16'hf227;
  rom[24570] = 16'he9e6;
  rom[24571] = 16'hea06;
  rom[24572] = 16'hf226;
  rom[24573] = 16'hea47;
  rom[24574] = 16'hd227;
  rom[24575] = 16'hdb2d;
  rom[24576] = 16'hff3c;
  rom[24577] = 16'hffff;
  rom[24578] = 16'hffff;
  rom[24579] = 16'hffff;
  rom[24580] = 16'hffff;
  rom[24581] = 16'hffff;
  rom[24582] = 16'hffff;
  rom[24583] = 16'hffff;
  rom[24584] = 16'hffff;
  rom[24585] = 16'hffff;
  rom[24586] = 16'hffff;
  rom[24587] = 16'hffff;
  rom[24588] = 16'hffff;
  rom[24589] = 16'hffff;
  rom[24590] = 16'hffff;
  rom[24591] = 16'hffff;
  rom[24592] = 16'hffff;
  rom[24593] = 16'hffff;
  rom[24594] = 16'hffff;
  rom[24595] = 16'hffff;
  rom[24596] = 16'hffff;
  rom[24597] = 16'hffff;
  rom[24598] = 16'hffff;
  rom[24599] = 16'hffff;
  rom[24600] = 16'hffff;
  rom[24601] = 16'hffff;
  rom[24602] = 16'hffff;
  rom[24603] = 16'hffff;
  rom[24604] = 16'hffff;
  rom[24605] = 16'hffff;
  rom[24606] = 16'hffff;
  rom[24607] = 16'hffff;
  rom[24608] = 16'hffff;
  rom[24609] = 16'hff7c;
  rom[24610] = 16'hc34d;
  rom[24611] = 16'hba89;
  rom[24612] = 16'hd36d;
  rom[24613] = 16'hf595;
  rom[24614] = 16'hff5c;
  rom[24615] = 16'hff9d;
  rom[24616] = 16'hffde;
  rom[24617] = 16'hffdf;
  rom[24618] = 16'hffff;
  rom[24619] = 16'hffff;
  rom[24620] = 16'hffff;
  rom[24621] = 16'hffff;
  rom[24622] = 16'hffff;
  rom[24623] = 16'hffff;
  rom[24624] = 16'hffff;
  rom[24625] = 16'hffff;
  rom[24626] = 16'hffff;
  rom[24627] = 16'hffff;
  rom[24628] = 16'hffff;
  rom[24629] = 16'hffff;
  rom[24630] = 16'hffff;
  rom[24631] = 16'hffff;
  rom[24632] = 16'hffff;
  rom[24633] = 16'hffff;
  rom[24634] = 16'hffff;
  rom[24635] = 16'hffff;
  rom[24636] = 16'hffdf;
  rom[24637] = 16'hfffe;
  rom[24638] = 16'hffdd;
  rom[24639] = 16'hff9b;
  rom[24640] = 16'hff3a;
  rom[24641] = 16'hf5b5;
  rom[24642] = 16'hdbee;
  rom[24643] = 16'hcaa8;
  rom[24644] = 16'hda68;
  rom[24645] = 16'hda26;
  rom[24646] = 16'hea48;
  rom[24647] = 16'hf227;
  rom[24648] = 16'hf207;
  rom[24649] = 16'hea05;
  rom[24650] = 16'hea86;
  rom[24651] = 16'he245;
  rom[24652] = 16'hea46;
  rom[24653] = 16'hea67;
  rom[24654] = 16'he248;
  rom[24655] = 16'hda49;
  rom[24656] = 16'hc227;
  rom[24657] = 16'h99a3;
  rom[24658] = 16'h7941;
  rom[24659] = 16'h9ac4;
  rom[24660] = 16'hdd4b;
  rom[24661] = 16'hfe8d;
  rom[24662] = 16'hfeec;
  rom[24663] = 16'hfeea;
  rom[24664] = 16'hfeea;
  rom[24665] = 16'hf6ea;
  rom[24666] = 16'hf74c;
  rom[24667] = 16'hf72b;
  rom[24668] = 16'hff2a;
  rom[24669] = 16'hff09;
  rom[24670] = 16'hff29;
  rom[24671] = 16'hff28;
  rom[24672] = 16'hf729;
  rom[24673] = 16'hf708;
  rom[24674] = 16'hff4a;
  rom[24675] = 16'hff2a;
  rom[24676] = 16'hfeea;
  rom[24677] = 16'hfeca;
  rom[24678] = 16'hff0c;
  rom[24679] = 16'hfeeb;
  rom[24680] = 16'hf6ee;
  rom[24681] = 16'he66d;
  rom[24682] = 16'hce0d;
  rom[24683] = 16'ha4ea;
  rom[24684] = 16'h83a7;
  rom[24685] = 16'h7326;
  rom[24686] = 16'h83a9;
  rom[24687] = 16'ha510;
  rom[24688] = 16'hd657;
  rom[24689] = 16'hef3b;
  rom[24690] = 16'hffdd;
  rom[24691] = 16'hffbd;
  rom[24692] = 16'hffde;
  rom[24693] = 16'hfffe;
  rom[24694] = 16'hffff;
  rom[24695] = 16'hffff;
  rom[24696] = 16'hffff;
  rom[24697] = 16'hffff;
  rom[24698] = 16'hffff;
  rom[24699] = 16'hffde;
  rom[24700] = 16'hffff;
  rom[24701] = 16'hffde;
  rom[24702] = 16'hffdf;
  rom[24703] = 16'hff9d;
  rom[24704] = 16'hff5c;
  rom[24705] = 16'heeb8;
  rom[24706] = 16'hcdd4;
  rom[24707] = 16'h944c;
  rom[24708] = 16'h7b88;
  rom[24709] = 16'h7386;
  rom[24710] = 16'h9489;
  rom[24711] = 16'hb56a;
  rom[24712] = 16'hde6d;
  rom[24713] = 16'heeee;
  rom[24714] = 16'hf70d;
  rom[24715] = 16'hf6ea;
  rom[24716] = 16'hff4a;
  rom[24717] = 16'hff49;
  rom[24718] = 16'hff49;
  rom[24719] = 16'hf749;
  rom[24720] = 16'hff2a;
  rom[24721] = 16'hf70a;
  rom[24722] = 16'hff2b;
  rom[24723] = 16'hff0a;
  rom[24724] = 16'hff0a;
  rom[24725] = 16'hff29;
  rom[24726] = 16'hf709;
  rom[24727] = 16'hf70a;
  rom[24728] = 16'hff0f;
  rom[24729] = 16'h7261;
  rom[24730] = 16'h6181;
  rom[24731] = 16'h59a1;
  rom[24732] = 16'hbcc9;
  rom[24733] = 16'he6cd;
  rom[24734] = 16'hef2c;
  rom[24735] = 16'hf74b;
  rom[24736] = 16'hf729;
  rom[24737] = 16'hf70a;
  rom[24738] = 16'hff4a;
  rom[24739] = 16'hf70a;
  rom[24740] = 16'hff2a;
  rom[24741] = 16'hf729;
  rom[24742] = 16'hff29;
  rom[24743] = 16'hff28;
  rom[24744] = 16'hff29;
  rom[24745] = 16'hff28;
  rom[24746] = 16'hff49;
  rom[24747] = 16'hf708;
  rom[24748] = 16'hff09;
  rom[24749] = 16'hfee8;
  rom[24750] = 16'hff29;
  rom[24751] = 16'hff09;
  rom[24752] = 16'hff29;
  rom[24753] = 16'hf72a;
  rom[24754] = 16'hff4d;
  rom[24755] = 16'hf6ed;
  rom[24756] = 16'hee2d;
  rom[24757] = 16'h9b66;
  rom[24758] = 16'h69a1;
  rom[24759] = 16'h9a65;
  rom[24760] = 16'hcaa7;
  rom[24761] = 16'he288;
  rom[24762] = 16'hea07;
  rom[24763] = 16'hf207;
  rom[24764] = 16'hfa07;
  rom[24765] = 16'hf1e6;
  rom[24766] = 16'hf226;
  rom[24767] = 16'hea26;
  rom[24768] = 16'hf227;
  rom[24769] = 16'hf1e7;
  rom[24770] = 16'hf9e7;
  rom[24771] = 16'hf1e6;
  rom[24772] = 16'hfa07;
  rom[24773] = 16'hf227;
  rom[24774] = 16'hda28;
  rom[24775] = 16'he34e;
  rom[24776] = 16'hff3d;
  rom[24777] = 16'hffff;
  rom[24778] = 16'hffff;
  rom[24779] = 16'hffff;
  rom[24780] = 16'hffff;
  rom[24781] = 16'hffff;
  rom[24782] = 16'hffff;
  rom[24783] = 16'hffff;
  rom[24784] = 16'hffff;
  rom[24785] = 16'hffff;
  rom[24786] = 16'hffff;
  rom[24787] = 16'hffff;
  rom[24788] = 16'hffff;
  rom[24789] = 16'hffff;
  rom[24790] = 16'hffff;
  rom[24791] = 16'hffff;
  rom[24792] = 16'hffff;
  rom[24793] = 16'hffff;
  rom[24794] = 16'hffff;
  rom[24795] = 16'hffff;
  rom[24796] = 16'hffff;
  rom[24797] = 16'hffff;
  rom[24798] = 16'hffff;
  rom[24799] = 16'hffff;
  rom[24800] = 16'hffff;
  rom[24801] = 16'hffff;
  rom[24802] = 16'hffff;
  rom[24803] = 16'hffff;
  rom[24804] = 16'hffdf;
  rom[24805] = 16'hffff;
  rom[24806] = 16'hffff;
  rom[24807] = 16'hffff;
  rom[24808] = 16'hffde;
  rom[24809] = 16'hff1b;
  rom[24810] = 16'hc289;
  rom[24811] = 16'he269;
  rom[24812] = 16'hda49;
  rom[24813] = 16'hcaca;
  rom[24814] = 16'hf4d2;
  rom[24815] = 16'hfe79;
  rom[24816] = 16'hff5c;
  rom[24817] = 16'hffff;
  rom[24818] = 16'hffff;
  rom[24819] = 16'hffff;
  rom[24820] = 16'hffff;
  rom[24821] = 16'hffdf;
  rom[24822] = 16'hffff;
  rom[24823] = 16'hffff;
  rom[24824] = 16'hffff;
  rom[24825] = 16'hffff;
  rom[24826] = 16'hffff;
  rom[24827] = 16'hffff;
  rom[24828] = 16'hffff;
  rom[24829] = 16'hffff;
  rom[24830] = 16'hffff;
  rom[24831] = 16'hffff;
  rom[24832] = 16'hffff;
  rom[24833] = 16'hffff;
  rom[24834] = 16'hffde;
  rom[24835] = 16'hffff;
  rom[24836] = 16'hffbd;
  rom[24837] = 16'hff9c;
  rom[24838] = 16'hff1a;
  rom[24839] = 16'hfdb4;
  rom[24840] = 16'hd3cd;
  rom[24841] = 16'hc288;
  rom[24842] = 16'hda68;
  rom[24843] = 16'he268;
  rom[24844] = 16'hda26;
  rom[24845] = 16'hda06;
  rom[24846] = 16'hea47;
  rom[24847] = 16'hea07;
  rom[24848] = 16'hea06;
  rom[24849] = 16'hf206;
  rom[24850] = 16'hf206;
  rom[24851] = 16'hf226;
  rom[24852] = 16'he9e6;
  rom[24853] = 16'he1c6;
  rom[24854] = 16'hea28;
  rom[24855] = 16'hf289;
  rom[24856] = 16'hda47;
  rom[24857] = 16'hda87;
  rom[24858] = 16'hc286;
  rom[24859] = 16'h8961;
  rom[24860] = 16'h6920;
  rom[24861] = 16'ha305;
  rom[24862] = 16'he5cd;
  rom[24863] = 16'heecc;
  rom[24864] = 16'hf72b;
  rom[24865] = 16'hff4c;
  rom[24866] = 16'hef0a;
  rom[24867] = 16'hff2a;
  rom[24868] = 16'hf709;
  rom[24869] = 16'hf709;
  rom[24870] = 16'hf709;
  rom[24871] = 16'hff49;
  rom[24872] = 16'hf729;
  rom[24873] = 16'hff69;
  rom[24874] = 16'hf707;
  rom[24875] = 16'hf728;
  rom[24876] = 16'hff69;
  rom[24877] = 16'hff29;
  rom[24878] = 16'hf70a;
  rom[24879] = 16'hff4b;
  rom[24880] = 16'heec9;
  rom[24881] = 16'heeca;
  rom[24882] = 16'hf70c;
  rom[24883] = 16'hf72e;
  rom[24884] = 16'hf72f;
  rom[24885] = 16'hf710;
  rom[24886] = 16'hbd4a;
  rom[24887] = 16'h9c49;
  rom[24888] = 16'h5a42;
  rom[24889] = 16'h49e3;
  rom[24890] = 16'h6ac6;
  rom[24891] = 16'h93eb;
  rom[24892] = 16'hac8e;
  rom[24893] = 16'hacb1;
  rom[24894] = 16'hb4f2;
  rom[24895] = 16'hc575;
  rom[24896] = 16'hde37;
  rom[24897] = 16'hee99;
  rom[24898] = 16'he5f6;
  rom[24899] = 16'hd574;
  rom[24900] = 16'hbcb1;
  rom[24901] = 16'hb42f;
  rom[24902] = 16'ha40d;
  rom[24903] = 16'h82e8;
  rom[24904] = 16'h5a03;
  rom[24905] = 16'h51e1;
  rom[24906] = 16'h7344;
  rom[24907] = 16'hb52b;
  rom[24908] = 16'hd66e;
  rom[24909] = 16'he6ee;
  rom[24910] = 16'heeed;
  rom[24911] = 16'hff2d;
  rom[24912] = 16'hff8d;
  rom[24913] = 16'hff2b;
  rom[24914] = 16'hfeea;
  rom[24915] = 16'hff4a;
  rom[24916] = 16'hf6e7;
  rom[24917] = 16'heee7;
  rom[24918] = 16'hf728;
  rom[24919] = 16'hf729;
  rom[24920] = 16'hf709;
  rom[24921] = 16'hff29;
  rom[24922] = 16'hff09;
  rom[24923] = 16'hff29;
  rom[24924] = 16'hef09;
  rom[24925] = 16'hf728;
  rom[24926] = 16'hf729;
  rom[24927] = 16'hff4d;
  rom[24928] = 16'he5eb;
  rom[24929] = 16'h71a0;
  rom[24930] = 16'ha286;
  rom[24931] = 16'h91a4;
  rom[24932] = 16'h6920;
  rom[24933] = 16'h9b87;
  rom[24934] = 16'he66e;
  rom[24935] = 16'hf70c;
  rom[24936] = 16'hff8b;
  rom[24937] = 16'hf70a;
  rom[24938] = 16'hf72a;
  rom[24939] = 16'hf709;
  rom[24940] = 16'hef29;
  rom[24941] = 16'hf749;
  rom[24942] = 16'hf709;
  rom[24943] = 16'hff2a;
  rom[24944] = 16'hf6e8;
  rom[24945] = 16'hff28;
  rom[24946] = 16'hf707;
  rom[24947] = 16'hff29;
  rom[24948] = 16'hf72a;
  rom[24949] = 16'hf709;
  rom[24950] = 16'hf709;
  rom[24951] = 16'hff49;
  rom[24952] = 16'hf728;
  rom[24953] = 16'hff49;
  rom[24954] = 16'hf709;
  rom[24955] = 16'hf70a;
  rom[24956] = 16'hf6ca;
  rom[24957] = 16'hff4e;
  rom[24958] = 16'hb4c7;
  rom[24959] = 16'h6160;
  rom[24960] = 16'h91c3;
  rom[24961] = 16'hc267;
  rom[24962] = 16'hd267;
  rom[24963] = 16'hea06;
  rom[24964] = 16'hfa07;
  rom[24965] = 16'hf9e7;
  rom[24966] = 16'hf207;
  rom[24967] = 16'hf227;
  rom[24968] = 16'he9e6;
  rom[24969] = 16'hfa27;
  rom[24970] = 16'hf1e6;
  rom[24971] = 16'hf207;
  rom[24972] = 16'hea26;
  rom[24973] = 16'hea48;
  rom[24974] = 16'hd227;
  rom[24975] = 16'he3cf;
  rom[24976] = 16'hff5d;
  rom[24977] = 16'hffff;
  rom[24978] = 16'hffff;
  rom[24979] = 16'hffff;
  rom[24980] = 16'hffff;
  rom[24981] = 16'hffff;
  rom[24982] = 16'hffff;
  rom[24983] = 16'hffff;
  rom[24984] = 16'hffff;
  rom[24985] = 16'hffff;
  rom[24986] = 16'hffff;
  rom[24987] = 16'hffff;
  rom[24988] = 16'hffff;
  rom[24989] = 16'hffff;
  rom[24990] = 16'hffff;
  rom[24991] = 16'hffff;
  rom[24992] = 16'hffff;
  rom[24993] = 16'hffff;
  rom[24994] = 16'hffff;
  rom[24995] = 16'hffff;
  rom[24996] = 16'hffff;
  rom[24997] = 16'hffff;
  rom[24998] = 16'hffff;
  rom[24999] = 16'hffff;
  rom[25000] = 16'hffff;
  rom[25001] = 16'hffff;
  rom[25002] = 16'hffff;
  rom[25003] = 16'hffff;
  rom[25004] = 16'hffff;
  rom[25005] = 16'hffff;
  rom[25006] = 16'hffff;
  rom[25007] = 16'hffff;
  rom[25008] = 16'hffde;
  rom[25009] = 16'hff1a;
  rom[25010] = 16'hd2a9;
  rom[25011] = 16'hea08;
  rom[25012] = 16'hf228;
  rom[25013] = 16'hda07;
  rom[25014] = 16'hd289;
  rom[25015] = 16'hdbad;
  rom[25016] = 16'hf554;
  rom[25017] = 16'hfeb9;
  rom[25018] = 16'hff9d;
  rom[25019] = 16'hffbe;
  rom[25020] = 16'hffff;
  rom[25021] = 16'hffff;
  rom[25022] = 16'hffff;
  rom[25023] = 16'hffff;
  rom[25024] = 16'hffff;
  rom[25025] = 16'hffff;
  rom[25026] = 16'hffff;
  rom[25027] = 16'hffff;
  rom[25028] = 16'hffff;
  rom[25029] = 16'hffff;
  rom[25030] = 16'hffff;
  rom[25031] = 16'hfffe;
  rom[25032] = 16'hffff;
  rom[25033] = 16'hffbd;
  rom[25034] = 16'hff9d;
  rom[25035] = 16'hff1b;
  rom[25036] = 16'hfe58;
  rom[25037] = 16'he4b1;
  rom[25038] = 16'hdbad;
  rom[25039] = 16'hd2c9;
  rom[25040] = 16'hda68;
  rom[25041] = 16'he227;
  rom[25042] = 16'hea07;
  rom[25043] = 16'hea06;
  rom[25044] = 16'hf248;
  rom[25045] = 16'hea48;
  rom[25046] = 16'hea07;
  rom[25047] = 16'hf227;
  rom[25048] = 16'hf207;
  rom[25049] = 16'hf206;
  rom[25050] = 16'hf1e7;
  rom[25051] = 16'hf1e6;
  rom[25052] = 16'hf206;
  rom[25053] = 16'hf227;
  rom[25054] = 16'hea07;
  rom[25055] = 16'he206;
  rom[25056] = 16'hea47;
  rom[25057] = 16'he226;
  rom[25058] = 16'he287;
  rom[25059] = 16'hca87;
  rom[25060] = 16'hb225;
  rom[25061] = 16'h8942;
  rom[25062] = 16'h79a2;
  rom[25063] = 16'h9b44;
  rom[25064] = 16'hcd67;
  rom[25065] = 16'heecd;
  rom[25066] = 16'hff0b;
  rom[25067] = 16'hff09;
  rom[25068] = 16'hff2a;
  rom[25069] = 16'hff29;
  rom[25070] = 16'hff2a;
  rom[25071] = 16'hf729;
  rom[25072] = 16'hff49;
  rom[25073] = 16'hf728;
  rom[25074] = 16'hff48;
  rom[25075] = 16'hff48;
  rom[25076] = 16'hf708;
  rom[25077] = 16'hf729;
  rom[25078] = 16'hff4a;
  rom[25079] = 16'hff09;
  rom[25080] = 16'hff29;
  rom[25081] = 16'hff29;
  rom[25082] = 16'hff0a;
  rom[25083] = 16'hff0a;
  rom[25084] = 16'hff0b;
  rom[25085] = 16'hf70c;
  rom[25086] = 16'hff0f;
  rom[25087] = 16'hfed0;
  rom[25088] = 16'hfeb1;
  rom[25089] = 16'hee10;
  rom[25090] = 16'he58f;
  rom[25091] = 16'hdd0d;
  rom[25092] = 16'hc44c;
  rom[25093] = 16'h9ac7;
  rom[25094] = 16'h81e6;
  rom[25095] = 16'h79e5;
  rom[25096] = 16'h8245;
  rom[25097] = 16'h8a65;
  rom[25098] = 16'h8a25;
  rom[25099] = 16'h79a4;
  rom[25100] = 16'h89c5;
  rom[25101] = 16'h9a26;
  rom[25102] = 16'haa47;
  rom[25103] = 16'hb348;
  rom[25104] = 16'hdd2d;
  rom[25105] = 16'hf690;
  rom[25106] = 16'hf710;
  rom[25107] = 16'hef6e;
  rom[25108] = 16'hf74d;
  rom[25109] = 16'hef2b;
  rom[25110] = 16'hff4b;
  rom[25111] = 16'hef09;
  rom[25112] = 16'hf709;
  rom[25113] = 16'hff09;
  rom[25114] = 16'hff0a;
  rom[25115] = 16'hf6e8;
  rom[25116] = 16'hff29;
  rom[25117] = 16'hff49;
  rom[25118] = 16'hff4a;
  rom[25119] = 16'hff29;
  rom[25120] = 16'hff2a;
  rom[25121] = 16'hff29;
  rom[25122] = 16'hff29;
  rom[25123] = 16'hff28;
  rom[25124] = 16'hf729;
  rom[25125] = 16'hf749;
  rom[25126] = 16'hff4a;
  rom[25127] = 16'hf6eb;
  rom[25128] = 16'hdd8b;
  rom[25129] = 16'h79a0;
  rom[25130] = 16'hba47;
  rom[25131] = 16'hca88;
  rom[25132] = 16'hb267;
  rom[25133] = 16'h7161;
  rom[25134] = 16'h8ae4;
  rom[25135] = 16'hd5ca;
  rom[25136] = 16'hf70c;
  rom[25137] = 16'hf72b;
  rom[25138] = 16'hf72a;
  rom[25139] = 16'hf729;
  rom[25140] = 16'hf74a;
  rom[25141] = 16'hef29;
  rom[25142] = 16'hff2a;
  rom[25143] = 16'hf709;
  rom[25144] = 16'hff29;
  rom[25145] = 16'hff08;
  rom[25146] = 16'hff49;
  rom[25147] = 16'hf709;
  rom[25148] = 16'hf72a;
  rom[25149] = 16'hff4a;
  rom[25150] = 16'hf709;
  rom[25151] = 16'hf708;
  rom[25152] = 16'hff49;
  rom[25153] = 16'hf728;
  rom[25154] = 16'hff4a;
  rom[25155] = 16'hff09;
  rom[25156] = 16'hff0a;
  rom[25157] = 16'hf72b;
  rom[25158] = 16'hf70c;
  rom[25159] = 16'hcd08;
  rom[25160] = 16'h8a43;
  rom[25161] = 16'h89a3;
  rom[25162] = 16'hcac8;
  rom[25163] = 16'hda67;
  rom[25164] = 16'hf227;
  rom[25165] = 16'hf207;
  rom[25166] = 16'hf227;
  rom[25167] = 16'he227;
  rom[25168] = 16'hea47;
  rom[25169] = 16'hea06;
  rom[25170] = 16'hf227;
  rom[25171] = 16'hea07;
  rom[25172] = 16'hea27;
  rom[25173] = 16'he227;
  rom[25174] = 16'hda89;
  rom[25175] = 16'hec2f;
  rom[25176] = 16'hff7d;
  rom[25177] = 16'hffff;
  rom[25178] = 16'hffff;
  rom[25179] = 16'hffff;
  rom[25180] = 16'hffff;
  rom[25181] = 16'hffff;
  rom[25182] = 16'hffff;
  rom[25183] = 16'hffff;
  rom[25184] = 16'hffff;
  rom[25185] = 16'hffff;
  rom[25186] = 16'hffff;
  rom[25187] = 16'hffff;
  rom[25188] = 16'hffff;
  rom[25189] = 16'hffff;
  rom[25190] = 16'hffff;
  rom[25191] = 16'hffff;
  rom[25192] = 16'hffff;
  rom[25193] = 16'hffff;
  rom[25194] = 16'hffff;
  rom[25195] = 16'hffff;
  rom[25196] = 16'hffff;
  rom[25197] = 16'hffff;
  rom[25198] = 16'hffff;
  rom[25199] = 16'hffff;
  rom[25200] = 16'hffff;
  rom[25201] = 16'hffff;
  rom[25202] = 16'hffff;
  rom[25203] = 16'hffff;
  rom[25204] = 16'hffff;
  rom[25205] = 16'hffff;
  rom[25206] = 16'hffff;
  rom[25207] = 16'hffff;
  rom[25208] = 16'hffde;
  rom[25209] = 16'hfeda;
  rom[25210] = 16'hd2a9;
  rom[25211] = 16'hea07;
  rom[25212] = 16'hea06;
  rom[25213] = 16'hea06;
  rom[25214] = 16'hda47;
  rom[25215] = 16'hda88;
  rom[25216] = 16'hcaa9;
  rom[25217] = 16'hd3ad;
  rom[25218] = 16'he4f2;
  rom[25219] = 16'hf5d5;
  rom[25220] = 16'hfef9;
  rom[25221] = 16'hff5a;
  rom[25222] = 16'hff9c;
  rom[25223] = 16'hffbd;
  rom[25224] = 16'hffbd;
  rom[25225] = 16'hffbe;
  rom[25226] = 16'hffde;
  rom[25227] = 16'hffbe;
  rom[25228] = 16'hff9d;
  rom[25229] = 16'hff7d;
  rom[25230] = 16'hff3b;
  rom[25231] = 16'hfefa;
  rom[25232] = 16'hfe98;
  rom[25233] = 16'hfdf7;
  rom[25234] = 16'hdcd1;
  rom[25235] = 16'hcb8d;
  rom[25236] = 16'hc2ca;
  rom[25237] = 16'hd269;
  rom[25238] = 16'he249;
  rom[25239] = 16'hea28;
  rom[25240] = 16'hea08;
  rom[25241] = 16'hfa48;
  rom[25242] = 16'he9e6;
  rom[25243] = 16'hea27;
  rom[25244] = 16'hea27;
  rom[25245] = 16'hea07;
  rom[25246] = 16'hea27;
  rom[25247] = 16'hea26;
  rom[25248] = 16'hf206;
  rom[25249] = 16'hf207;
  rom[25250] = 16'hf227;
  rom[25251] = 16'hf206;
  rom[25252] = 16'hf207;
  rom[25253] = 16'hf206;
  rom[25254] = 16'he1e6;
  rom[25255] = 16'hea27;
  rom[25256] = 16'hea27;
  rom[25257] = 16'hea27;
  rom[25258] = 16'he226;
  rom[25259] = 16'hd226;
  rom[25260] = 16'hd267;
  rom[25261] = 16'hd289;
  rom[25262] = 16'hb226;
  rom[25263] = 16'h89e2;
  rom[25264] = 16'h6180;
  rom[25265] = 16'h9b86;
  rom[25266] = 16'hf6cb;
  rom[25267] = 16'hff09;
  rom[25268] = 16'hf708;
  rom[25269] = 16'hff29;
  rom[25270] = 16'hf709;
  rom[25271] = 16'hf729;
  rom[25272] = 16'hff29;
  rom[25273] = 16'hff48;
  rom[25274] = 16'hf728;
  rom[25275] = 16'hf728;
  rom[25276] = 16'hff69;
  rom[25277] = 16'hf729;
  rom[25278] = 16'hf708;
  rom[25279] = 16'hff28;
  rom[25280] = 16'hff27;
  rom[25281] = 16'hf6c6;
  rom[25282] = 16'hff08;
  rom[25283] = 16'hff09;
  rom[25284] = 16'hf72a;
  rom[25285] = 16'hff6d;
  rom[25286] = 16'hf6ab;
  rom[25287] = 16'hfe6c;
  rom[25288] = 16'hfdcb;
  rom[25289] = 16'hf4ea;
  rom[25290] = 16'hf4ca;
  rom[25291] = 16'hdbe8;
  rom[25292] = 16'hd388;
  rom[25293] = 16'hba86;
  rom[25294] = 16'hc2c8;
  rom[25295] = 16'hcae8;
  rom[25296] = 16'hcb48;
  rom[25297] = 16'hecad;
  rom[25298] = 16'hc327;
  rom[25299] = 16'hc2e7;
  rom[25300] = 16'hcaa7;
  rom[25301] = 16'hca47;
  rom[25302] = 16'hd225;
  rom[25303] = 16'hd2c6;
  rom[25304] = 16'hdbe7;
  rom[25305] = 16'hfe8e;
  rom[25306] = 16'hf70c;
  rom[25307] = 16'he70a;
  rom[25308] = 16'he709;
  rom[25309] = 16'hf729;
  rom[25310] = 16'hf708;
  rom[25311] = 16'hff49;
  rom[25312] = 16'hf708;
  rom[25313] = 16'hff2a;
  rom[25314] = 16'hff0a;
  rom[25315] = 16'hff49;
  rom[25316] = 16'hff29;
  rom[25317] = 16'hff29;
  rom[25318] = 16'hf708;
  rom[25319] = 16'hff29;
  rom[25320] = 16'hff09;
  rom[25321] = 16'hff29;
  rom[25322] = 16'hf709;
  rom[25323] = 16'hff28;
  rom[25324] = 16'hf729;
  rom[25325] = 16'hf708;
  rom[25326] = 16'hf789;
  rom[25327] = 16'hf72c;
  rom[25328] = 16'hb4a7;
  rom[25329] = 16'h6941;
  rom[25330] = 16'hca88;
  rom[25331] = 16'he2a8;
  rom[25332] = 16'hd267;
  rom[25333] = 16'hc2a8;
  rom[25334] = 16'h7960;
  rom[25335] = 16'h7a21;
  rom[25336] = 16'hcd69;
  rom[25337] = 16'hfeed;
  rom[25338] = 16'hf72b;
  rom[25339] = 16'hf70a;
  rom[25340] = 16'hef09;
  rom[25341] = 16'hff8b;
  rom[25342] = 16'heee8;
  rom[25343] = 16'hff49;
  rom[25344] = 16'hff08;
  rom[25345] = 16'hff29;
  rom[25346] = 16'hf709;
  rom[25347] = 16'hf729;
  rom[25348] = 16'hf709;
  rom[25349] = 16'hff2a;
  rom[25350] = 16'hf729;
  rom[25351] = 16'hff29;
  rom[25352] = 16'hf728;
  rom[25353] = 16'hff48;
  rom[25354] = 16'hf708;
  rom[25355] = 16'hff6a;
  rom[25356] = 16'hf709;
  rom[25357] = 16'hff2b;
  rom[25358] = 16'hf72a;
  rom[25359] = 16'hf6cb;
  rom[25360] = 16'he5cc;
  rom[25361] = 16'h8222;
  rom[25362] = 16'h89c2;
  rom[25363] = 16'hcaa7;
  rom[25364] = 16'he267;
  rom[25365] = 16'hea26;
  rom[25366] = 16'he226;
  rom[25367] = 16'he247;
  rom[25368] = 16'he226;
  rom[25369] = 16'hea27;
  rom[25370] = 16'hea26;
  rom[25371] = 16'hea06;
  rom[25372] = 16'hea27;
  rom[25373] = 16'hea27;
  rom[25374] = 16'hd268;
  rom[25375] = 16'hecd1;
  rom[25376] = 16'hff7c;
  rom[25377] = 16'hffff;
  rom[25378] = 16'hffff;
  rom[25379] = 16'hffff;
  rom[25380] = 16'hffff;
  rom[25381] = 16'hffff;
  rom[25382] = 16'hffff;
  rom[25383] = 16'hffff;
  rom[25384] = 16'hffff;
  rom[25385] = 16'hffff;
  rom[25386] = 16'hffff;
  rom[25387] = 16'hffff;
  rom[25388] = 16'hffff;
  rom[25389] = 16'hffff;
  rom[25390] = 16'hffff;
  rom[25391] = 16'hffff;
  rom[25392] = 16'hffff;
  rom[25393] = 16'hffff;
  rom[25394] = 16'hffff;
  rom[25395] = 16'hffff;
  rom[25396] = 16'hffff;
  rom[25397] = 16'hffff;
  rom[25398] = 16'hffff;
  rom[25399] = 16'hffff;
  rom[25400] = 16'hffff;
  rom[25401] = 16'hffff;
  rom[25402] = 16'hffff;
  rom[25403] = 16'hffff;
  rom[25404] = 16'hffff;
  rom[25405] = 16'hffff;
  rom[25406] = 16'hffff;
  rom[25407] = 16'hffff;
  rom[25408] = 16'hffff;
  rom[25409] = 16'hfe78;
  rom[25410] = 16'hd2a9;
  rom[25411] = 16'hea26;
  rom[25412] = 16'hf246;
  rom[25413] = 16'hea05;
  rom[25414] = 16'hf247;
  rom[25415] = 16'hea27;
  rom[25416] = 16'he228;
  rom[25417] = 16'hda48;
  rom[25418] = 16'hd289;
  rom[25419] = 16'hcaea;
  rom[25420] = 16'he3cd;
  rom[25421] = 16'hecb0;
  rom[25422] = 16'hf512;
  rom[25423] = 16'hf595;
  rom[25424] = 16'hfdd7;
  rom[25425] = 16'hf5d6;
  rom[25426] = 16'hfdd7;
  rom[25427] = 16'hf5d6;
  rom[25428] = 16'hf5b5;
  rom[25429] = 16'hf574;
  rom[25430] = 16'hf4f2;
  rom[25431] = 16'he40e;
  rom[25432] = 16'hdb6c;
  rom[25433] = 16'hdaea;
  rom[25434] = 16'hd2a9;
  rom[25435] = 16'hd268;
  rom[25436] = 16'he268;
  rom[25437] = 16'he207;
  rom[25438] = 16'hf247;
  rom[25439] = 16'hea07;
  rom[25440] = 16'hf207;
  rom[25441] = 16'hea07;
  rom[25442] = 16'hf227;
  rom[25443] = 16'hea07;
  rom[25444] = 16'hf228;
  rom[25445] = 16'hf227;
  rom[25446] = 16'hea07;
  rom[25447] = 16'hea27;
  rom[25448] = 16'hf227;
  rom[25449] = 16'hf206;
  rom[25450] = 16'hf206;
  rom[25451] = 16'hf206;
  rom[25452] = 16'hf227;
  rom[25453] = 16'hf207;
  rom[25454] = 16'hf227;
  rom[25455] = 16'hea27;
  rom[25456] = 16'hea27;
  rom[25457] = 16'hf227;
  rom[25458] = 16'hea27;
  rom[25459] = 16'he246;
  rom[25460] = 16'hea47;
  rom[25461] = 16'hea49;
  rom[25462] = 16'hda4a;
  rom[25463] = 16'hc288;
  rom[25464] = 16'h89e2;
  rom[25465] = 16'h92e4;
  rom[25466] = 16'hfeee;
  rom[25467] = 16'hf74a;
  rom[25468] = 16'hff29;
  rom[25469] = 16'hff29;
  rom[25470] = 16'hff2a;
  rom[25471] = 16'hff29;
  rom[25472] = 16'hff2a;
  rom[25473] = 16'hff28;
  rom[25474] = 16'hf729;
  rom[25475] = 16'hff28;
  rom[25476] = 16'hf708;
  rom[25477] = 16'hf729;
  rom[25478] = 16'hff49;
  rom[25479] = 16'hff28;
  rom[25480] = 16'hff08;
  rom[25481] = 16'hff29;
  rom[25482] = 16'hff29;
  rom[25483] = 16'hf709;
  rom[25484] = 16'hff2a;
  rom[25485] = 16'hfeea;
  rom[25486] = 16'hfe8b;
  rom[25487] = 16'hd4a4;
  rom[25488] = 16'hcb82;
  rom[25489] = 16'hc2e1;
  rom[25490] = 16'hd2c3;
  rom[25491] = 16'hd284;
  rom[25492] = 16'hda65;
  rom[25493] = 16'hda46;
  rom[25494] = 16'hda88;
  rom[25495] = 16'hba45;
  rom[25496] = 16'hdbe9;
  rom[25497] = 16'hfd6f;
  rom[25498] = 16'hf4cd;
  rom[25499] = 16'hcac7;
  rom[25500] = 16'hd267;
  rom[25501] = 16'hea47;
  rom[25502] = 16'hf227;
  rom[25503] = 16'hea45;
  rom[25504] = 16'hdac3;
  rom[25505] = 16'hfd69;
  rom[25506] = 16'hfeec;
  rom[25507] = 16'hf729;
  rom[25508] = 16'hff49;
  rom[25509] = 16'hff08;
  rom[25510] = 16'hff29;
  rom[25511] = 16'hf749;
  rom[25512] = 16'hf728;
  rom[25513] = 16'hff2a;
  rom[25514] = 16'hff0a;
  rom[25515] = 16'hff08;
  rom[25516] = 16'hff29;
  rom[25517] = 16'hf728;
  rom[25518] = 16'hff29;
  rom[25519] = 16'hff29;
  rom[25520] = 16'hff2a;
  rom[25521] = 16'hff29;
  rom[25522] = 16'hff29;
  rom[25523] = 16'hff28;
  rom[25524] = 16'hff49;
  rom[25525] = 16'hf728;
  rom[25526] = 16'hf749;
  rom[25527] = 16'hef2b;
  rom[25528] = 16'h9c47;
  rom[25529] = 16'h7182;
  rom[25530] = 16'hd248;
  rom[25531] = 16'he1e5;
  rom[25532] = 16'hea27;
  rom[25533] = 16'he288;
  rom[25534] = 16'hba66;
  rom[25535] = 16'h89e2;
  rom[25536] = 16'h79e1;
  rom[25537] = 16'hcd29;
  rom[25538] = 16'hff0d;
  rom[25539] = 16'hf72a;
  rom[25540] = 16'hff4a;
  rom[25541] = 16'hf6c9;
  rom[25542] = 16'hff4a;
  rom[25543] = 16'hf708;
  rom[25544] = 16'hff29;
  rom[25545] = 16'hff09;
  rom[25546] = 16'hff2a;
  rom[25547] = 16'hff29;
  rom[25548] = 16'hff4a;
  rom[25549] = 16'hf709;
  rom[25550] = 16'hff2a;
  rom[25551] = 16'hf729;
  rom[25552] = 16'hff49;
  rom[25553] = 16'hf728;
  rom[25554] = 16'hff49;
  rom[25555] = 16'hf708;
  rom[25556] = 16'hff29;
  rom[25557] = 16'hf709;
  rom[25558] = 16'hff29;
  rom[25559] = 16'hf6e9;
  rom[25560] = 16'hf6ed;
  rom[25561] = 16'hc54a;
  rom[25562] = 16'h79e1;
  rom[25563] = 16'ha204;
  rom[25564] = 16'hd246;
  rom[25565] = 16'he246;
  rom[25566] = 16'he227;
  rom[25567] = 16'he248;
  rom[25568] = 16'he268;
  rom[25569] = 16'hea27;
  rom[25570] = 16'hf227;
  rom[25571] = 16'hea06;
  rom[25572] = 16'hf227;
  rom[25573] = 16'hea07;
  rom[25574] = 16'hdaa9;
  rom[25575] = 16'hed53;
  rom[25576] = 16'hfffe;
  rom[25577] = 16'hffff;
  rom[25578] = 16'hffff;
  rom[25579] = 16'hffff;
  rom[25580] = 16'hffff;
  rom[25581] = 16'hffff;
  rom[25582] = 16'hffff;
  rom[25583] = 16'hffff;
  rom[25584] = 16'hffff;
  rom[25585] = 16'hffff;
  rom[25586] = 16'hffff;
  rom[25587] = 16'hffff;
  rom[25588] = 16'hffff;
  rom[25589] = 16'hffff;
  rom[25590] = 16'hffff;
  rom[25591] = 16'hffff;
  rom[25592] = 16'hffff;
  rom[25593] = 16'hffff;
  rom[25594] = 16'hffff;
  rom[25595] = 16'hffff;
  rom[25596] = 16'hffff;
  rom[25597] = 16'hffff;
  rom[25598] = 16'hffff;
  rom[25599] = 16'hffff;
  rom[25600] = 16'hffff;
  rom[25601] = 16'hffff;
  rom[25602] = 16'hffff;
  rom[25603] = 16'hffff;
  rom[25604] = 16'hffff;
  rom[25605] = 16'hffff;
  rom[25606] = 16'hffff;
  rom[25607] = 16'hffff;
  rom[25608] = 16'hffde;
  rom[25609] = 16'hf617;
  rom[25610] = 16'hd269;
  rom[25611] = 16'hea47;
  rom[25612] = 16'he1e5;
  rom[25613] = 16'hea26;
  rom[25614] = 16'hea07;
  rom[25615] = 16'hf207;
  rom[25616] = 16'hea07;
  rom[25617] = 16'hf208;
  rom[25618] = 16'hea08;
  rom[25619] = 16'he248;
  rom[25620] = 16'hda27;
  rom[25621] = 16'hd207;
  rom[25622] = 16'hda69;
  rom[25623] = 16'hdaaa;
  rom[25624] = 16'hdaaa;
  rom[25625] = 16'hdacb;
  rom[25626] = 16'hd2ca;
  rom[25627] = 16'hd2cb;
  rom[25628] = 16'hcaca;
  rom[25629] = 16'hd2a9;
  rom[25630] = 16'hca68;
  rom[25631] = 16'hda88;
  rom[25632] = 16'he268;
  rom[25633] = 16'hea47;
  rom[25634] = 16'hea47;
  rom[25635] = 16'hea27;
  rom[25636] = 16'he227;
  rom[25637] = 16'hea47;
  rom[25638] = 16'hea47;
  rom[25639] = 16'hea26;
  rom[25640] = 16'hea06;
  rom[25641] = 16'hea27;
  rom[25642] = 16'hf227;
  rom[25643] = 16'hf227;
  rom[25644] = 16'hea07;
  rom[25645] = 16'hea07;
  rom[25646] = 16'hea07;
  rom[25647] = 16'hea07;
  rom[25648] = 16'he9e6;
  rom[25649] = 16'hea06;
  rom[25650] = 16'hea27;
  rom[25651] = 16'hf226;
  rom[25652] = 16'he9e6;
  rom[25653] = 16'hea27;
  rom[25654] = 16'hea27;
  rom[25655] = 16'hf227;
  rom[25656] = 16'hea27;
  rom[25657] = 16'hea27;
  rom[25658] = 16'hea47;
  rom[25659] = 16'hea46;
  rom[25660] = 16'he224;
  rom[25661] = 16'hf207;
  rom[25662] = 16'hda48;
  rom[25663] = 16'hd2a9;
  rom[25664] = 16'haa65;
  rom[25665] = 16'h7224;
  rom[25666] = 16'he68c;
  rom[25667] = 16'hef0a;
  rom[25668] = 16'hf728;
  rom[25669] = 16'hff28;
  rom[25670] = 16'hff09;
  rom[25671] = 16'hff29;
  rom[25672] = 16'hf709;
  rom[25673] = 16'hf709;
  rom[25674] = 16'hff49;
  rom[25675] = 16'hff29;
  rom[25676] = 16'hf748;
  rom[25677] = 16'hf729;
  rom[25678] = 16'hf708;
  rom[25679] = 16'hf729;
  rom[25680] = 16'hef09;
  rom[25681] = 16'hf729;
  rom[25682] = 16'hf729;
  rom[25683] = 16'hf6e9;
  rom[25684] = 16'hff2a;
  rom[25685] = 16'hf6aa;
  rom[25686] = 16'hbc42;
  rom[25687] = 16'hcc43;
  rom[25688] = 16'hdc86;
  rom[25689] = 16'he426;
  rom[25690] = 16'hdb45;
  rom[25691] = 16'hd264;
  rom[25692] = 16'hda66;
  rom[25693] = 16'hd226;
  rom[25694] = 16'hca26;
  rom[25695] = 16'hc286;
  rom[25696] = 16'hd3e9;
  rom[25697] = 16'hed0c;
  rom[25698] = 16'heced;
  rom[25699] = 16'hdb89;
  rom[25700] = 16'hd2c8;
  rom[25701] = 16'he248;
  rom[25702] = 16'hd9e7;
  rom[25703] = 16'hda06;
  rom[25704] = 16'hdac5;
  rom[25705] = 16'hdba4;
  rom[25706] = 16'hf5c9;
  rom[25707] = 16'hfeca;
  rom[25708] = 16'hfec8;
  rom[25709] = 16'hfee8;
  rom[25710] = 16'hff09;
  rom[25711] = 16'hf729;
  rom[25712] = 16'hef8a;
  rom[25713] = 16'hff2a;
  rom[25714] = 16'hff09;
  rom[25715] = 16'hff29;
  rom[25716] = 16'hf728;
  rom[25717] = 16'hff29;
  rom[25718] = 16'hf708;
  rom[25719] = 16'hff29;
  rom[25720] = 16'hf709;
  rom[25721] = 16'hff29;
  rom[25722] = 16'hff09;
  rom[25723] = 16'hff28;
  rom[25724] = 16'hf708;
  rom[25725] = 16'hff28;
  rom[25726] = 16'he6e8;
  rom[25727] = 16'hf74c;
  rom[25728] = 16'h8ba5;
  rom[25729] = 16'h79a3;
  rom[25730] = 16'hd227;
  rom[25731] = 16'hfa06;
  rom[25732] = 16'hf9c5;
  rom[25733] = 16'he9c6;
  rom[25734] = 16'hd227;
  rom[25735] = 16'hc2a7;
  rom[25736] = 16'h9a24;
  rom[25737] = 16'h8242;
  rom[25738] = 16'hcd49;
  rom[25739] = 16'hf70d;
  rom[25740] = 16'hf72a;
  rom[25741] = 16'hff4a;
  rom[25742] = 16'hf708;
  rom[25743] = 16'hff49;
  rom[25744] = 16'hf709;
  rom[25745] = 16'hff49;
  rom[25746] = 16'hff09;
  rom[25747] = 16'hf709;
  rom[25748] = 16'hf708;
  rom[25749] = 16'hff49;
  rom[25750] = 16'hff09;
  rom[25751] = 16'hff29;
  rom[25752] = 16'hf728;
  rom[25753] = 16'hff29;
  rom[25754] = 16'hf708;
  rom[25755] = 16'hff49;
  rom[25756] = 16'hf708;
  rom[25757] = 16'hff29;
  rom[25758] = 16'hff07;
  rom[25759] = 16'hff28;
  rom[25760] = 16'hf70a;
  rom[25761] = 16'hf6ee;
  rom[25762] = 16'hc4e9;
  rom[25763] = 16'h81c1;
  rom[25764] = 16'hba65;
  rom[25765] = 16'hda67;
  rom[25766] = 16'he228;
  rom[25767] = 16'he207;
  rom[25768] = 16'he226;
  rom[25769] = 16'hea26;
  rom[25770] = 16'hea26;
  rom[25771] = 16'hfa47;
  rom[25772] = 16'he9e6;
  rom[25773] = 16'hea07;
  rom[25774] = 16'hdac9;
  rom[25775] = 16'hf5f5;
  rom[25776] = 16'hffdd;
  rom[25777] = 16'hffff;
  rom[25778] = 16'hffff;
  rom[25779] = 16'hffff;
  rom[25780] = 16'hffff;
  rom[25781] = 16'hffff;
  rom[25782] = 16'hffff;
  rom[25783] = 16'hffff;
  rom[25784] = 16'hffff;
  rom[25785] = 16'hffff;
  rom[25786] = 16'hffff;
  rom[25787] = 16'hffff;
  rom[25788] = 16'hffff;
  rom[25789] = 16'hffff;
  rom[25790] = 16'hffff;
  rom[25791] = 16'hffff;
  rom[25792] = 16'hffff;
  rom[25793] = 16'hffff;
  rom[25794] = 16'hffff;
  rom[25795] = 16'hffff;
  rom[25796] = 16'hffff;
  rom[25797] = 16'hffff;
  rom[25798] = 16'hffff;
  rom[25799] = 16'hffff;
  rom[25800] = 16'hffff;
  rom[25801] = 16'hffff;
  rom[25802] = 16'hffff;
  rom[25803] = 16'hffff;
  rom[25804] = 16'hffff;
  rom[25805] = 16'hffff;
  rom[25806] = 16'hffff;
  rom[25807] = 16'hffff;
  rom[25808] = 16'hffff;
  rom[25809] = 16'hf616;
  rom[25810] = 16'hda89;
  rom[25811] = 16'hea48;
  rom[25812] = 16'he9c6;
  rom[25813] = 16'hf227;
  rom[25814] = 16'hf207;
  rom[25815] = 16'hf227;
  rom[25816] = 16'hfa28;
  rom[25817] = 16'hf228;
  rom[25818] = 16'hf208;
  rom[25819] = 16'he9c7;
  rom[25820] = 16'hf229;
  rom[25821] = 16'hf208;
  rom[25822] = 16'hf208;
  rom[25823] = 16'hea28;
  rom[25824] = 16'hea28;
  rom[25825] = 16'he207;
  rom[25826] = 16'hea48;
  rom[25827] = 16'hea48;
  rom[25828] = 16'he248;
  rom[25829] = 16'he247;
  rom[25830] = 16'hea67;
  rom[25831] = 16'hea47;
  rom[25832] = 16'hea26;
  rom[25833] = 16'he9e6;
  rom[25834] = 16'hf207;
  rom[25835] = 16'hf206;
  rom[25836] = 16'hf247;
  rom[25837] = 16'he226;
  rom[25838] = 16'hea47;
  rom[25839] = 16'hea26;
  rom[25840] = 16'hea26;
  rom[25841] = 16'hf227;
  rom[25842] = 16'hf227;
  rom[25843] = 16'hea27;
  rom[25844] = 16'hea27;
  rom[25845] = 16'hea27;
  rom[25846] = 16'hf227;
  rom[25847] = 16'hea27;
  rom[25848] = 16'hf247;
  rom[25849] = 16'hea26;
  rom[25850] = 16'hea27;
  rom[25851] = 16'hea26;
  rom[25852] = 16'hf247;
  rom[25853] = 16'hea26;
  rom[25854] = 16'hea27;
  rom[25855] = 16'hea07;
  rom[25856] = 16'hea27;
  rom[25857] = 16'hf227;
  rom[25858] = 16'hea07;
  rom[25859] = 16'hea45;
  rom[25860] = 16'hf245;
  rom[25861] = 16'hea05;
  rom[25862] = 16'he228;
  rom[25863] = 16'hd267;
  rom[25864] = 16'hbaa6;
  rom[25865] = 16'h69a2;
  rom[25866] = 16'hde4c;
  rom[25867] = 16'hef2a;
  rom[25868] = 16'hff49;
  rom[25869] = 16'hff29;
  rom[25870] = 16'hff2a;
  rom[25871] = 16'hff29;
  rom[25872] = 16'hff2a;
  rom[25873] = 16'hff29;
  rom[25874] = 16'hff09;
  rom[25875] = 16'hff29;
  rom[25876] = 16'hf729;
  rom[25877] = 16'hf728;
  rom[25878] = 16'hff49;
  rom[25879] = 16'hf729;
  rom[25880] = 16'hf72a;
  rom[25881] = 16'hff4b;
  rom[25882] = 16'hf72a;
  rom[25883] = 16'hff2a;
  rom[25884] = 16'hff2a;
  rom[25885] = 16'hee27;
  rom[25886] = 16'he586;
  rom[25887] = 16'hfe0a;
  rom[25888] = 16'hfe8e;
  rom[25889] = 16'hfe0d;
  rom[25890] = 16'hf4ec;
  rom[25891] = 16'he3aa;
  rom[25892] = 16'hb9e5;
  rom[25893] = 16'ha923;
  rom[25894] = 16'ha102;
  rom[25895] = 16'h9941;
  rom[25896] = 16'h8982;
  rom[25897] = 16'h8a02;
  rom[25898] = 16'h9a43;
  rom[25899] = 16'ha203;
  rom[25900] = 16'ha963;
  rom[25901] = 16'hb9a6;
  rom[25902] = 16'hda4a;
  rom[25903] = 16'hda89;
  rom[25904] = 16'hd2c7;
  rom[25905] = 16'hbaa3;
  rom[25906] = 16'hcbe4;
  rom[25907] = 16'he545;
  rom[25908] = 16'hfea9;
  rom[25909] = 16'hfec8;
  rom[25910] = 16'hff2a;
  rom[25911] = 16'hf74a;
  rom[25912] = 16'he72a;
  rom[25913] = 16'hff09;
  rom[25914] = 16'hff0a;
  rom[25915] = 16'hff29;
  rom[25916] = 16'hff29;
  rom[25917] = 16'hff28;
  rom[25918] = 16'hff49;
  rom[25919] = 16'hff29;
  rom[25920] = 16'hff2a;
  rom[25921] = 16'hff29;
  rom[25922] = 16'hff29;
  rom[25923] = 16'hff28;
  rom[25924] = 16'hff29;
  rom[25925] = 16'hff49;
  rom[25926] = 16'hf709;
  rom[25927] = 16'heecc;
  rom[25928] = 16'h7b24;
  rom[25929] = 16'h9246;
  rom[25930] = 16'he248;
  rom[25931] = 16'hf9e5;
  rom[25932] = 16'hf9c5;
  rom[25933] = 16'hf9e8;
  rom[25934] = 16'hea09;
  rom[25935] = 16'hd227;
  rom[25936] = 16'hcaa7;
  rom[25937] = 16'h99c3;
  rom[25938] = 16'h8242;
  rom[25939] = 16'hcd49;
  rom[25940] = 16'heecb;
  rom[25941] = 16'hf729;
  rom[25942] = 16'hff49;
  rom[25943] = 16'hf728;
  rom[25944] = 16'hff49;
  rom[25945] = 16'hf6e8;
  rom[25946] = 16'hff4a;
  rom[25947] = 16'hff29;
  rom[25948] = 16'hff2a;
  rom[25949] = 16'hff29;
  rom[25950] = 16'hf72a;
  rom[25951] = 16'hff29;
  rom[25952] = 16'hff4a;
  rom[25953] = 16'hf728;
  rom[25954] = 16'hff4a;
  rom[25955] = 16'hff28;
  rom[25956] = 16'hff49;
  rom[25957] = 16'hff28;
  rom[25958] = 16'hff28;
  rom[25959] = 16'hf6e8;
  rom[25960] = 16'hff6b;
  rom[25961] = 16'heeeb;
  rom[25962] = 16'hff4f;
  rom[25963] = 16'hab84;
  rom[25964] = 16'h8960;
  rom[25965] = 16'hca46;
  rom[25966] = 16'he249;
  rom[25967] = 16'hea28;
  rom[25968] = 16'hea27;
  rom[25969] = 16'hea27;
  rom[25970] = 16'hea06;
  rom[25971] = 16'hf227;
  rom[25972] = 16'hf207;
  rom[25973] = 16'hf227;
  rom[25974] = 16'hdaeb;
  rom[25975] = 16'hf657;
  rom[25976] = 16'hfffe;
  rom[25977] = 16'hffff;
  rom[25978] = 16'hffff;
  rom[25979] = 16'hffff;
  rom[25980] = 16'hffff;
  rom[25981] = 16'hffff;
  rom[25982] = 16'hffff;
  rom[25983] = 16'hffff;
  rom[25984] = 16'hffff;
  rom[25985] = 16'hffff;
  rom[25986] = 16'hffff;
  rom[25987] = 16'hffff;
  rom[25988] = 16'hffff;
  rom[25989] = 16'hffff;
  rom[25990] = 16'hffff;
  rom[25991] = 16'hffff;
  rom[25992] = 16'hffff;
  rom[25993] = 16'hffff;
  rom[25994] = 16'hffff;
  rom[25995] = 16'hffff;
  rom[25996] = 16'hffff;
  rom[25997] = 16'hffff;
  rom[25998] = 16'hffff;
  rom[25999] = 16'hffff;
  rom[26000] = 16'hfffe;
  rom[26001] = 16'hffff;
  rom[26002] = 16'hffff;
  rom[26003] = 16'hffff;
  rom[26004] = 16'hffff;
  rom[26005] = 16'hffff;
  rom[26006] = 16'hffff;
  rom[26007] = 16'hffff;
  rom[26008] = 16'hffde;
  rom[26009] = 16'hfe99;
  rom[26010] = 16'hd269;
  rom[26011] = 16'hea28;
  rom[26012] = 16'hf207;
  rom[26013] = 16'hf227;
  rom[26014] = 16'he9e7;
  rom[26015] = 16'hf1e7;
  rom[26016] = 16'hea07;
  rom[26017] = 16'hea07;
  rom[26018] = 16'he9e6;
  rom[26019] = 16'hea08;
  rom[26020] = 16'hf207;
  rom[26021] = 16'hf228;
  rom[26022] = 16'hea07;
  rom[26023] = 16'hf226;
  rom[26024] = 16'hea26;
  rom[26025] = 16'hf206;
  rom[26026] = 16'hea06;
  rom[26027] = 16'hf227;
  rom[26028] = 16'hea27;
  rom[26029] = 16'hea27;
  rom[26030] = 16'he206;
  rom[26031] = 16'he226;
  rom[26032] = 16'hea26;
  rom[26033] = 16'hf227;
  rom[26034] = 16'hea06;
  rom[26035] = 16'hf207;
  rom[26036] = 16'hf206;
  rom[26037] = 16'hf226;
  rom[26038] = 16'hea06;
  rom[26039] = 16'hf227;
  rom[26040] = 16'hf206;
  rom[26041] = 16'hf206;
  rom[26042] = 16'hea06;
  rom[26043] = 16'hea26;
  rom[26044] = 16'hea26;
  rom[26045] = 16'hea07;
  rom[26046] = 16'hea06;
  rom[26047] = 16'hea06;
  rom[26048] = 16'hea26;
  rom[26049] = 16'hea26;
  rom[26050] = 16'he226;
  rom[26051] = 16'hea26;
  rom[26052] = 16'hea26;
  rom[26053] = 16'hea26;
  rom[26054] = 16'he206;
  rom[26055] = 16'hf207;
  rom[26056] = 16'hea07;
  rom[26057] = 16'hf207;
  rom[26058] = 16'hea06;
  rom[26059] = 16'hea26;
  rom[26060] = 16'hea25;
  rom[26061] = 16'hf226;
  rom[26062] = 16'he227;
  rom[26063] = 16'hda67;
  rom[26064] = 16'hc285;
  rom[26065] = 16'h71a1;
  rom[26066] = 16'hd5ea;
  rom[26067] = 16'hef2b;
  rom[26068] = 16'hf708;
  rom[26069] = 16'hff29;
  rom[26070] = 16'hf709;
  rom[26071] = 16'hff29;
  rom[26072] = 16'hff29;
  rom[26073] = 16'hff29;
  rom[26074] = 16'hf709;
  rom[26075] = 16'hff29;
  rom[26076] = 16'hff09;
  rom[26077] = 16'hff28;
  rom[26078] = 16'hf728;
  rom[26079] = 16'hf748;
  rom[26080] = 16'hf728;
  rom[26081] = 16'hf729;
  rom[26082] = 16'hf729;
  rom[26083] = 16'hff4a;
  rom[26084] = 16'hff28;
  rom[26085] = 16'hf6a7;
  rom[26086] = 16'hfec9;
  rom[26087] = 16'hfecc;
  rom[26088] = 16'hfeae;
  rom[26089] = 16'hedee;
  rom[26090] = 16'hc429;
  rom[26091] = 16'h89c4;
  rom[26092] = 16'h9963;
  rom[26093] = 16'hb184;
  rom[26094] = 16'hc1e4;
  rom[26095] = 16'hc225;
  rom[26096] = 16'hc246;
  rom[26097] = 16'hb225;
  rom[26098] = 16'hb244;
  rom[26099] = 16'hba24;
  rom[26100] = 16'ha963;
  rom[26101] = 16'ha103;
  rom[26102] = 16'h90c3;
  rom[26103] = 16'hb227;
  rom[26104] = 16'hdbab;
  rom[26105] = 16'hec8b;
  rom[26106] = 16'he4e8;
  rom[26107] = 16'hed87;
  rom[26108] = 16'hee26;
  rom[26109] = 16'hff08;
  rom[26110] = 16'hf748;
  rom[26111] = 16'hf749;
  rom[26112] = 16'hef28;
  rom[26113] = 16'hff09;
  rom[26114] = 16'hff09;
  rom[26115] = 16'hff29;
  rom[26116] = 16'hf708;
  rom[26117] = 16'hff48;
  rom[26118] = 16'hf708;
  rom[26119] = 16'hff28;
  rom[26120] = 16'hff09;
  rom[26121] = 16'hff29;
  rom[26122] = 16'hf708;
  rom[26123] = 16'hff28;
  rom[26124] = 16'hff08;
  rom[26125] = 16'hff29;
  rom[26126] = 16'heec9;
  rom[26127] = 16'he66b;
  rom[26128] = 16'h7262;
  rom[26129] = 16'ha267;
  rom[26130] = 16'hda47;
  rom[26131] = 16'hf225;
  rom[26132] = 16'hf9e5;
  rom[26133] = 16'hf9e7;
  rom[26134] = 16'hf1e8;
  rom[26135] = 16'he227;
  rom[26136] = 16'hda66;
  rom[26137] = 16'hd267;
  rom[26138] = 16'h91c3;
  rom[26139] = 16'h8242;
  rom[26140] = 16'hd5aa;
  rom[26141] = 16'hf70b;
  rom[26142] = 16'hf729;
  rom[26143] = 16'hff29;
  rom[26144] = 16'hf708;
  rom[26145] = 16'hff4a;
  rom[26146] = 16'hf708;
  rom[26147] = 16'hff49;
  rom[26148] = 16'hf708;
  rom[26149] = 16'hff29;
  rom[26150] = 16'hf708;
  rom[26151] = 16'hff29;
  rom[26152] = 16'hff09;
  rom[26153] = 16'hff29;
  rom[26154] = 16'hf709;
  rom[26155] = 16'hff28;
  rom[26156] = 16'hff08;
  rom[26157] = 16'hff28;
  rom[26158] = 16'hff09;
  rom[26159] = 16'hff4a;
  rom[26160] = 16'hf709;
  rom[26161] = 16'hff4a;
  rom[26162] = 16'heec8;
  rom[26163] = 16'hedea;
  rom[26164] = 16'h8a21;
  rom[26165] = 16'ha1c4;
  rom[26166] = 16'hca48;
  rom[26167] = 16'he228;
  rom[26168] = 16'hea06;
  rom[26169] = 16'hf227;
  rom[26170] = 16'he9e6;
  rom[26171] = 16'hf226;
  rom[26172] = 16'hf206;
  rom[26173] = 16'hea28;
  rom[26174] = 16'hdb6c;
  rom[26175] = 16'hfef9;
  rom[26176] = 16'hfffe;
  rom[26177] = 16'hffff;
  rom[26178] = 16'hffff;
  rom[26179] = 16'hffff;
  rom[26180] = 16'hffff;
  rom[26181] = 16'hffff;
  rom[26182] = 16'hffff;
  rom[26183] = 16'hffff;
  rom[26184] = 16'hffff;
  rom[26185] = 16'hffff;
  rom[26186] = 16'hffff;
  rom[26187] = 16'hffff;
  rom[26188] = 16'hffff;
  rom[26189] = 16'hffff;
  rom[26190] = 16'hffff;
  rom[26191] = 16'hffff;
  rom[26192] = 16'hffff;
  rom[26193] = 16'hffff;
  rom[26194] = 16'hffff;
  rom[26195] = 16'hffff;
  rom[26196] = 16'hffff;
  rom[26197] = 16'hffff;
  rom[26198] = 16'hffff;
  rom[26199] = 16'hffff;
  rom[26200] = 16'hffff;
  rom[26201] = 16'hffff;
  rom[26202] = 16'hffff;
  rom[26203] = 16'hffff;
  rom[26204] = 16'hffff;
  rom[26205] = 16'hffff;
  rom[26206] = 16'hffff;
  rom[26207] = 16'hffff;
  rom[26208] = 16'hffff;
  rom[26209] = 16'hfefa;
  rom[26210] = 16'hd2ca;
  rom[26211] = 16'he207;
  rom[26212] = 16'hf268;
  rom[26213] = 16'hf206;
  rom[26214] = 16'hf247;
  rom[26215] = 16'hf206;
  rom[26216] = 16'hf248;
  rom[26217] = 16'hf227;
  rom[26218] = 16'hf247;
  rom[26219] = 16'hea27;
  rom[26220] = 16'hea27;
  rom[26221] = 16'he206;
  rom[26222] = 16'he226;
  rom[26223] = 16'hea26;
  rom[26224] = 16'hea47;
  rom[26225] = 16'hea26;
  rom[26226] = 16'hf225;
  rom[26227] = 16'hf206;
  rom[26228] = 16'hf227;
  rom[26229] = 16'hf206;
  rom[26230] = 16'hea26;
  rom[26231] = 16'hea06;
  rom[26232] = 16'hea27;
  rom[26233] = 16'hea27;
  rom[26234] = 16'hea47;
  rom[26235] = 16'hea27;
  rom[26236] = 16'hf208;
  rom[26237] = 16'hf1e7;
  rom[26238] = 16'hf1e6;
  rom[26239] = 16'hf1e6;
  rom[26240] = 16'hf227;
  rom[26241] = 16'hf206;
  rom[26242] = 16'hf226;
  rom[26243] = 16'hea26;
  rom[26244] = 16'hf227;
  rom[26245] = 16'hf206;
  rom[26246] = 16'hf226;
  rom[26247] = 16'hea06;
  rom[26248] = 16'hea27;
  rom[26249] = 16'hea26;
  rom[26250] = 16'hea46;
  rom[26251] = 16'hea26;
  rom[26252] = 16'hea27;
  rom[26253] = 16'hea06;
  rom[26254] = 16'hea26;
  rom[26255] = 16'hf206;
  rom[26256] = 16'hf227;
  rom[26257] = 16'hf207;
  rom[26258] = 16'hfa29;
  rom[26259] = 16'hea07;
  rom[26260] = 16'hf227;
  rom[26261] = 16'hf207;
  rom[26262] = 16'he227;
  rom[26263] = 16'he247;
  rom[26264] = 16'hd2c7;
  rom[26265] = 16'h7961;
  rom[26266] = 16'hddab;
  rom[26267] = 16'hf72b;
  rom[26268] = 16'hf72a;
  rom[26269] = 16'hff29;
  rom[26270] = 16'hff49;
  rom[26271] = 16'hff28;
  rom[26272] = 16'hff2a;
  rom[26273] = 16'hff29;
  rom[26274] = 16'hff2a;
  rom[26275] = 16'hff29;
  rom[26276] = 16'hff2a;
  rom[26277] = 16'hff28;
  rom[26278] = 16'hff29;
  rom[26279] = 16'hff28;
  rom[26280] = 16'hff49;
  rom[26281] = 16'hff08;
  rom[26282] = 16'hff09;
  rom[26283] = 16'hff08;
  rom[26284] = 16'hff29;
  rom[26285] = 16'hff4a;
  rom[26286] = 16'hf6eb;
  rom[26287] = 16'hfeee;
  rom[26288] = 16'he56c;
  rom[26289] = 16'h8a42;
  rom[26290] = 16'h7940;
  rom[26291] = 16'hc308;
  rom[26292] = 16'hcaa8;
  rom[26293] = 16'hda87;
  rom[26294] = 16'he265;
  rom[26295] = 16'he266;
  rom[26296] = 16'hda28;
  rom[26297] = 16'hdaa9;
  rom[26298] = 16'hd266;
  rom[26299] = 16'hd265;
  rom[26300] = 16'hd245;
  rom[26301] = 16'hd267;
  rom[26302] = 16'hba26;
  rom[26303] = 16'h9121;
  rom[26304] = 16'hb286;
  rom[26305] = 16'hfd90;
  rom[26306] = 16'hfe90;
  rom[26307] = 16'hfeed;
  rom[26308] = 16'hff4b;
  rom[26309] = 16'hff49;
  rom[26310] = 16'hf748;
  rom[26311] = 16'hf728;
  rom[26312] = 16'hff29;
  rom[26313] = 16'hff09;
  rom[26314] = 16'hff2a;
  rom[26315] = 16'hff29;
  rom[26316] = 16'hff29;
  rom[26317] = 16'hff28;
  rom[26318] = 16'hff29;
  rom[26319] = 16'hff28;
  rom[26320] = 16'hff2a;
  rom[26321] = 16'hff28;
  rom[26322] = 16'hff29;
  rom[26323] = 16'hff28;
  rom[26324] = 16'hff29;
  rom[26325] = 16'hff29;
  rom[26326] = 16'hf6c9;
  rom[26327] = 16'hde0b;
  rom[26328] = 16'h71c1;
  rom[26329] = 16'haa67;
  rom[26330] = 16'hda68;
  rom[26331] = 16'hf225;
  rom[26332] = 16'hfa26;
  rom[26333] = 16'hf1c6;
  rom[26334] = 16'hf1c8;
  rom[26335] = 16'hf207;
  rom[26336] = 16'hea27;
  rom[26337] = 16'hda27;
  rom[26338] = 16'hd2a8;
  rom[26339] = 16'h89a2;
  rom[26340] = 16'h8283;
  rom[26341] = 16'hde2c;
  rom[26342] = 16'hff0c;
  rom[26343] = 16'hff4a;
  rom[26344] = 16'hff29;
  rom[26345] = 16'hf708;
  rom[26346] = 16'hff4a;
  rom[26347] = 16'hf709;
  rom[26348] = 16'hff2a;
  rom[26349] = 16'hff29;
  rom[26350] = 16'hf709;
  rom[26351] = 16'hff29;
  rom[26352] = 16'hff2a;
  rom[26353] = 16'hff29;
  rom[26354] = 16'hff2a;
  rom[26355] = 16'hff28;
  rom[26356] = 16'hff29;
  rom[26357] = 16'hff28;
  rom[26358] = 16'hf72a;
  rom[26359] = 16'hff4b;
  rom[26360] = 16'hf70a;
  rom[26361] = 16'hf728;
  rom[26362] = 16'heee7;
  rom[26363] = 16'hff2c;
  rom[26364] = 16'hc4c8;
  rom[26365] = 16'h7981;
  rom[26366] = 16'hc267;
  rom[26367] = 16'he247;
  rom[26368] = 16'hf227;
  rom[26369] = 16'hf206;
  rom[26370] = 16'hf226;
  rom[26371] = 16'hf1e5;
  rom[26372] = 16'hfa07;
  rom[26373] = 16'hd227;
  rom[26374] = 16'hdc0f;
  rom[26375] = 16'hff7c;
  rom[26376] = 16'hffff;
  rom[26377] = 16'hffff;
  rom[26378] = 16'hffff;
  rom[26379] = 16'hffff;
  rom[26380] = 16'hffff;
  rom[26381] = 16'hffff;
  rom[26382] = 16'hffff;
  rom[26383] = 16'hffff;
  rom[26384] = 16'hffff;
  rom[26385] = 16'hffff;
  rom[26386] = 16'hffff;
  rom[26387] = 16'hffff;
  rom[26388] = 16'hffff;
  rom[26389] = 16'hffff;
  rom[26390] = 16'hffff;
  rom[26391] = 16'hffff;
  rom[26392] = 16'hffff;
  rom[26393] = 16'hffff;
  rom[26394] = 16'hffff;
  rom[26395] = 16'hffff;
  rom[26396] = 16'hffff;
  rom[26397] = 16'hffff;
  rom[26398] = 16'hffff;
  rom[26399] = 16'hffff;
  rom[26400] = 16'hffff;
  rom[26401] = 16'hffff;
  rom[26402] = 16'hffff;
  rom[26403] = 16'hffff;
  rom[26404] = 16'hffff;
  rom[26405] = 16'hffff;
  rom[26406] = 16'hffff;
  rom[26407] = 16'hffff;
  rom[26408] = 16'hffde;
  rom[26409] = 16'hfefa;
  rom[26410] = 16'hd2ca;
  rom[26411] = 16'he228;
  rom[26412] = 16'hf267;
  rom[26413] = 16'hea26;
  rom[26414] = 16'hea46;
  rom[26415] = 16'hea26;
  rom[26416] = 16'hea06;
  rom[26417] = 16'hf226;
  rom[26418] = 16'hf206;
  rom[26419] = 16'hf226;
  rom[26420] = 16'hea26;
  rom[26421] = 16'hea26;
  rom[26422] = 16'hea26;
  rom[26423] = 16'hea46;
  rom[26424] = 16'hea26;
  rom[26425] = 16'hf226;
  rom[26426] = 16'hf206;
  rom[26427] = 16'hf226;
  rom[26428] = 16'hea06;
  rom[26429] = 16'hf227;
  rom[26430] = 16'hf206;
  rom[26431] = 16'hf207;
  rom[26432] = 16'hea07;
  rom[26433] = 16'hea07;
  rom[26434] = 16'hea06;
  rom[26435] = 16'hea27;
  rom[26436] = 16'hea07;
  rom[26437] = 16'hf207;
  rom[26438] = 16'hf207;
  rom[26439] = 16'hf227;
  rom[26440] = 16'hea06;
  rom[26441] = 16'hea26;
  rom[26442] = 16'hea26;
  rom[26443] = 16'hea26;
  rom[26444] = 16'hea06;
  rom[26445] = 16'hf206;
  rom[26446] = 16'hea06;
  rom[26447] = 16'hea06;
  rom[26448] = 16'hea06;
  rom[26449] = 16'hea06;
  rom[26450] = 16'hea06;
  rom[26451] = 16'hf206;
  rom[26452] = 16'hea06;
  rom[26453] = 16'hea06;
  rom[26454] = 16'hea06;
  rom[26455] = 16'hf226;
  rom[26456] = 16'hea06;
  rom[26457] = 16'hf206;
  rom[26458] = 16'hf1e8;
  rom[26459] = 16'hea08;
  rom[26460] = 16'he9e7;
  rom[26461] = 16'hf208;
  rom[26462] = 16'hea08;
  rom[26463] = 16'he248;
  rom[26464] = 16'hd266;
  rom[26465] = 16'h8141;
  rom[26466] = 16'hd529;
  rom[26467] = 16'hff2b;
  rom[26468] = 16'hf709;
  rom[26469] = 16'hf729;
  rom[26470] = 16'hff29;
  rom[26471] = 16'hff28;
  rom[26472] = 16'hf728;
  rom[26473] = 16'hff29;
  rom[26474] = 16'hff09;
  rom[26475] = 16'hff29;
  rom[26476] = 16'hf709;
  rom[26477] = 16'hff28;
  rom[26478] = 16'hff08;
  rom[26479] = 16'hff09;
  rom[26480] = 16'hff49;
  rom[26481] = 16'hfec7;
  rom[26482] = 16'hff08;
  rom[26483] = 16'hff09;
  rom[26484] = 16'hff4a;
  rom[26485] = 16'hf70b;
  rom[26486] = 16'hfecc;
  rom[26487] = 16'hc487;
  rom[26488] = 16'h9241;
  rom[26489] = 16'h9a03;
  rom[26490] = 16'hc2c6;
  rom[26491] = 16'hc284;
  rom[26492] = 16'hcaa4;
  rom[26493] = 16'hd2c4;
  rom[26494] = 16'hdaa3;
  rom[26495] = 16'hda84;
  rom[26496] = 16'hd265;
  rom[26497] = 16'hdaa6;
  rom[26498] = 16'hca64;
  rom[26499] = 16'hd2a3;
  rom[26500] = 16'hd2e2;
  rom[26501] = 16'hcac3;
  rom[26502] = 16'hc284;
  rom[26503] = 16'hc285;
  rom[26504] = 16'h99a2;
  rom[26505] = 16'h9203;
  rom[26506] = 16'hd4ca;
  rom[26507] = 16'hff10;
  rom[26508] = 16'heeeb;
  rom[26509] = 16'hf74a;
  rom[26510] = 16'hef28;
  rom[26511] = 16'hff48;
  rom[26512] = 16'hf6e7;
  rom[26513] = 16'hff4a;
  rom[26514] = 16'hf6e9;
  rom[26515] = 16'hff29;
  rom[26516] = 16'hf708;
  rom[26517] = 16'hff28;
  rom[26518] = 16'hff28;
  rom[26519] = 16'hff28;
  rom[26520] = 16'hf709;
  rom[26521] = 16'hff28;
  rom[26522] = 16'hff08;
  rom[26523] = 16'hff28;
  rom[26524] = 16'hf708;
  rom[26525] = 16'hff29;
  rom[26526] = 16'hfeea;
  rom[26527] = 16'hddcb;
  rom[26528] = 16'h7180;
  rom[26529] = 16'hc288;
  rom[26530] = 16'hda27;
  rom[26531] = 16'hf227;
  rom[26532] = 16'hea25;
  rom[26533] = 16'hf226;
  rom[26534] = 16'hf1e7;
  rom[26535] = 16'hf207;
  rom[26536] = 16'hea06;
  rom[26537] = 16'hf248;
  rom[26538] = 16'hd227;
  rom[26539] = 16'hba67;
  rom[26540] = 16'h7962;
  rom[26541] = 16'h8ac2;
  rom[26542] = 16'he60b;
  rom[26543] = 16'hff4c;
  rom[26544] = 16'hf6e8;
  rom[26545] = 16'hff4a;
  rom[26546] = 16'hf709;
  rom[26547] = 16'hff0a;
  rom[26548] = 16'hf729;
  rom[26549] = 16'hf729;
  rom[26550] = 16'hff48;
  rom[26551] = 16'hff28;
  rom[26552] = 16'hf708;
  rom[26553] = 16'hff29;
  rom[26554] = 16'hff09;
  rom[26555] = 16'hff29;
  rom[26556] = 16'hf708;
  rom[26557] = 16'hff29;
  rom[26558] = 16'hf70a;
  rom[26559] = 16'hf72b;
  rom[26560] = 16'hf709;
  rom[26561] = 16'hf728;
  rom[26562] = 16'hf748;
  rom[26563] = 16'hf72a;
  rom[26564] = 16'hde2c;
  rom[26565] = 16'h8283;
  rom[26566] = 16'ha1e4;
  rom[26567] = 16'hda68;
  rom[26568] = 16'he226;
  rom[26569] = 16'hf227;
  rom[26570] = 16'hea26;
  rom[26571] = 16'he9e5;
  rom[26572] = 16'hea27;
  rom[26573] = 16'hd289;
  rom[26574] = 16'hdcb2;
  rom[26575] = 16'hff9e;
  rom[26576] = 16'hffff;
  rom[26577] = 16'hffff;
  rom[26578] = 16'hffff;
  rom[26579] = 16'hffff;
  rom[26580] = 16'hffff;
  rom[26581] = 16'hffff;
  rom[26582] = 16'hffff;
  rom[26583] = 16'hffff;
  rom[26584] = 16'hffff;
  rom[26585] = 16'hffff;
  rom[26586] = 16'hffff;
  rom[26587] = 16'hffff;
  rom[26588] = 16'hffff;
  rom[26589] = 16'hffff;
  rom[26590] = 16'hffff;
  rom[26591] = 16'hffff;
  rom[26592] = 16'hffff;
  rom[26593] = 16'hffff;
  rom[26594] = 16'hffff;
  rom[26595] = 16'hffff;
  rom[26596] = 16'hffff;
  rom[26597] = 16'hffff;
  rom[26598] = 16'hffff;
  rom[26599] = 16'hffff;
  rom[26600] = 16'hffff;
  rom[26601] = 16'hffff;
  rom[26602] = 16'hffff;
  rom[26603] = 16'hffff;
  rom[26604] = 16'hffff;
  rom[26605] = 16'hffff;
  rom[26606] = 16'hffff;
  rom[26607] = 16'hffff;
  rom[26608] = 16'hffff;
  rom[26609] = 16'hff3b;
  rom[26610] = 16'hd2aa;
  rom[26611] = 16'hda27;
  rom[26612] = 16'hea87;
  rom[26613] = 16'hea26;
  rom[26614] = 16'hf247;
  rom[26615] = 16'hea06;
  rom[26616] = 16'hf226;
  rom[26617] = 16'hf226;
  rom[26618] = 16'hf226;
  rom[26619] = 16'hf206;
  rom[26620] = 16'hf226;
  rom[26621] = 16'hf206;
  rom[26622] = 16'hf206;
  rom[26623] = 16'hea06;
  rom[26624] = 16'hf226;
  rom[26625] = 16'hea06;
  rom[26626] = 16'hea27;
  rom[26627] = 16'hea06;
  rom[26628] = 16'hea26;
  rom[26629] = 16'hea06;
  rom[26630] = 16'hf228;
  rom[26631] = 16'hf207;
  rom[26632] = 16'hf207;
  rom[26633] = 16'hf1e7;
  rom[26634] = 16'hf227;
  rom[26635] = 16'hf206;
  rom[26636] = 16'hf227;
  rom[26637] = 16'hea07;
  rom[26638] = 16'hea27;
  rom[26639] = 16'hea26;
  rom[26640] = 16'hea46;
  rom[26641] = 16'hea26;
  rom[26642] = 16'hea47;
  rom[26643] = 16'hea26;
  rom[26644] = 16'hf226;
  rom[26645] = 16'hea26;
  rom[26646] = 16'hea27;
  rom[26647] = 16'hea06;
  rom[26648] = 16'hf226;
  rom[26649] = 16'hf206;
  rom[26650] = 16'hf227;
  rom[26651] = 16'hf206;
  rom[26652] = 16'hf226;
  rom[26653] = 16'hea06;
  rom[26654] = 16'hea27;
  rom[26655] = 16'hea26;
  rom[26656] = 16'hf226;
  rom[26657] = 16'hf206;
  rom[26658] = 16'hf1e8;
  rom[26659] = 16'hea07;
  rom[26660] = 16'hea27;
  rom[26661] = 16'hea07;
  rom[26662] = 16'hea28;
  rom[26663] = 16'he227;
  rom[26664] = 16'hda67;
  rom[26665] = 16'h9182;
  rom[26666] = 16'hc487;
  rom[26667] = 16'hff2b;
  rom[26668] = 16'hff2b;
  rom[26669] = 16'hf729;
  rom[26670] = 16'hff29;
  rom[26671] = 16'hff28;
  rom[26672] = 16'hff49;
  rom[26673] = 16'hff28;
  rom[26674] = 16'hff29;
  rom[26675] = 16'hff29;
  rom[26676] = 16'hff2a;
  rom[26677] = 16'hff28;
  rom[26678] = 16'hff29;
  rom[26679] = 16'hff09;
  rom[26680] = 16'hff09;
  rom[26681] = 16'hfee8;
  rom[26682] = 16'hff6a;
  rom[26683] = 16'hf709;
  rom[26684] = 16'hf70c;
  rom[26685] = 16'hff0e;
  rom[26686] = 16'hd50a;
  rom[26687] = 16'h8200;
  rom[26688] = 16'haa43;
  rom[26689] = 16'hcac5;
  rom[26690] = 16'hcac4;
  rom[26691] = 16'hf407;
  rom[26692] = 16'hfd49;
  rom[26693] = 16'hfd68;
  rom[26694] = 16'hfd49;
  rom[26695] = 16'hfd09;
  rom[26696] = 16'hfd0b;
  rom[26697] = 16'hfceb;
  rom[26698] = 16'hfd2c;
  rom[26699] = 16'hfd69;
  rom[26700] = 16'hfd87;
  rom[26701] = 16'hfda8;
  rom[26702] = 16'hf487;
  rom[26703] = 16'hd2e4;
  rom[26704] = 16'hca85;
  rom[26705] = 16'haa03;
  rom[26706] = 16'h8a02;
  rom[26707] = 16'he5ac;
  rom[26708] = 16'hff4e;
  rom[26709] = 16'hef2a;
  rom[26710] = 16'hf709;
  rom[26711] = 16'hff29;
  rom[26712] = 16'hf6e9;
  rom[26713] = 16'hf729;
  rom[26714] = 16'hf729;
  rom[26715] = 16'hff29;
  rom[26716] = 16'hff29;
  rom[26717] = 16'hff28;
  rom[26718] = 16'hff29;
  rom[26719] = 16'hff28;
  rom[26720] = 16'hff2a;
  rom[26721] = 16'hff28;
  rom[26722] = 16'hff29;
  rom[26723] = 16'hff29;
  rom[26724] = 16'hff2a;
  rom[26725] = 16'hff29;
  rom[26726] = 16'hfeeb;
  rom[26727] = 16'hcd29;
  rom[26728] = 16'h89c1;
  rom[26729] = 16'hca66;
  rom[26730] = 16'hea48;
  rom[26731] = 16'hf1e7;
  rom[26732] = 16'hea46;
  rom[26733] = 16'he246;
  rom[26734] = 16'hf228;
  rom[26735] = 16'hf206;
  rom[26736] = 16'hfa27;
  rom[26737] = 16'he9e6;
  rom[26738] = 16'hea69;
  rom[26739] = 16'hda88;
  rom[26740] = 16'hb247;
  rom[26741] = 16'h8181;
  rom[26742] = 16'habc6;
  rom[26743] = 16'hfecd;
  rom[26744] = 16'hff2c;
  rom[26745] = 16'hf6e8;
  rom[26746] = 16'hff2a;
  rom[26747] = 16'hf70a;
  rom[26748] = 16'hf72a;
  rom[26749] = 16'hff28;
  rom[26750] = 16'hff49;
  rom[26751] = 16'hf708;
  rom[26752] = 16'hff29;
  rom[26753] = 16'hff28;
  rom[26754] = 16'hff29;
  rom[26755] = 16'hff29;
  rom[26756] = 16'hff29;
  rom[26757] = 16'hff29;
  rom[26758] = 16'hff2a;
  rom[26759] = 16'hf729;
  rom[26760] = 16'hff49;
  rom[26761] = 16'hf707;
  rom[26762] = 16'hf708;
  rom[26763] = 16'hf76b;
  rom[26764] = 16'heeed;
  rom[26765] = 16'ha3a5;
  rom[26766] = 16'h99c3;
  rom[26767] = 16'hd267;
  rom[26768] = 16'he247;
  rom[26769] = 16'hf247;
  rom[26770] = 16'hea06;
  rom[26771] = 16'hf247;
  rom[26772] = 16'he227;
  rom[26773] = 16'hc2ca;
  rom[26774] = 16'hfe7a;
  rom[26775] = 16'hffbf;
  rom[26776] = 16'hffff;
  rom[26777] = 16'hffff;
  rom[26778] = 16'hffff;
  rom[26779] = 16'hffff;
  rom[26780] = 16'hffff;
  rom[26781] = 16'hffff;
  rom[26782] = 16'hffff;
  rom[26783] = 16'hffff;
  rom[26784] = 16'hffff;
  rom[26785] = 16'hffff;
  rom[26786] = 16'hffff;
  rom[26787] = 16'hffff;
  rom[26788] = 16'hffff;
  rom[26789] = 16'hffff;
  rom[26790] = 16'hffff;
  rom[26791] = 16'hffff;
  rom[26792] = 16'hffff;
  rom[26793] = 16'hffff;
  rom[26794] = 16'hffff;
  rom[26795] = 16'hffff;
  rom[26796] = 16'hffff;
  rom[26797] = 16'hffff;
  rom[26798] = 16'hffff;
  rom[26799] = 16'hffff;
  rom[26800] = 16'hffff;
  rom[26801] = 16'hffff;
  rom[26802] = 16'hffff;
  rom[26803] = 16'hffff;
  rom[26804] = 16'hffff;
  rom[26805] = 16'hffff;
  rom[26806] = 16'hffff;
  rom[26807] = 16'hffff;
  rom[26808] = 16'hffff;
  rom[26809] = 16'hff9d;
  rom[26810] = 16'hcaaa;
  rom[26811] = 16'he248;
  rom[26812] = 16'hea06;
  rom[26813] = 16'hea27;
  rom[26814] = 16'he206;
  rom[26815] = 16'hea26;
  rom[26816] = 16'hea06;
  rom[26817] = 16'hf207;
  rom[26818] = 16'he9e6;
  rom[26819] = 16'hf1e6;
  rom[26820] = 16'hf9e6;
  rom[26821] = 16'hfa06;
  rom[26822] = 16'hf1e6;
  rom[26823] = 16'hf207;
  rom[26824] = 16'hf207;
  rom[26825] = 16'hf207;
  rom[26826] = 16'hea27;
  rom[26827] = 16'hea27;
  rom[26828] = 16'hea27;
  rom[26829] = 16'hea27;
  rom[26830] = 16'hea27;
  rom[26831] = 16'hf227;
  rom[26832] = 16'hf207;
  rom[26833] = 16'hfa07;
  rom[26834] = 16'hf1e6;
  rom[26835] = 16'hf206;
  rom[26836] = 16'hf206;
  rom[26837] = 16'hf227;
  rom[26838] = 16'he226;
  rom[26839] = 16'hea27;
  rom[26840] = 16'hea27;
  rom[26841] = 16'hea27;
  rom[26842] = 16'hea07;
  rom[26843] = 16'hea27;
  rom[26844] = 16'hea26;
  rom[26845] = 16'hea26;
  rom[26846] = 16'he226;
  rom[26847] = 16'hea26;
  rom[26848] = 16'hea06;
  rom[26849] = 16'hf207;
  rom[26850] = 16'hea06;
  rom[26851] = 16'hf206;
  rom[26852] = 16'hf206;
  rom[26853] = 16'hf226;
  rom[26854] = 16'hea26;
  rom[26855] = 16'hea26;
  rom[26856] = 16'hea26;
  rom[26857] = 16'hea26;
  rom[26858] = 16'hea07;
  rom[26859] = 16'hea26;
  rom[26860] = 16'hea25;
  rom[26861] = 16'hea25;
  rom[26862] = 16'he225;
  rom[26863] = 16'hea46;
  rom[26864] = 16'hda46;
  rom[26865] = 16'ha1e4;
  rom[26866] = 16'h9b63;
  rom[26867] = 16'hf72b;
  rom[26868] = 16'hf70b;
  rom[26869] = 16'hf709;
  rom[26870] = 16'hf729;
  rom[26871] = 16'hff28;
  rom[26872] = 16'hff28;
  rom[26873] = 16'hff28;
  rom[26874] = 16'hf708;
  rom[26875] = 16'hff29;
  rom[26876] = 16'hff09;
  rom[26877] = 16'hff28;
  rom[26878] = 16'hf708;
  rom[26879] = 16'hff29;
  rom[26880] = 16'hf728;
  rom[26881] = 16'hff89;
  rom[26882] = 16'hef27;
  rom[26883] = 16'hef49;
  rom[26884] = 16'heeec;
  rom[26885] = 16'hd56b;
  rom[26886] = 16'h79e0;
  rom[26887] = 16'haa84;
  rom[26888] = 16'hcb06;
  rom[26889] = 16'hcac4;
  rom[26890] = 16'hd3a3;
  rom[26891] = 16'hfe09;
  rom[26892] = 16'hfec8;
  rom[26893] = 16'hfee8;
  rom[26894] = 16'hfea8;
  rom[26895] = 16'hfe08;
  rom[26896] = 16'hfda7;
  rom[26897] = 16'hfd88;
  rom[26898] = 16'hfdc9;
  rom[26899] = 16'hfeea;
  rom[26900] = 16'hff05;
  rom[26901] = 16'hff27;
  rom[26902] = 16'hfda6;
  rom[26903] = 16'hd321;
  rom[26904] = 16'hd283;
  rom[26905] = 16'hd286;
  rom[26906] = 16'ha203;
  rom[26907] = 16'h8a20;
  rom[26908] = 16'he60b;
  rom[26909] = 16'hff6d;
  rom[26910] = 16'hf709;
  rom[26911] = 16'hff69;
  rom[26912] = 16'hf708;
  rom[26913] = 16'hff29;
  rom[26914] = 16'hf708;
  rom[26915] = 16'hff29;
  rom[26916] = 16'hf728;
  rom[26917] = 16'hff48;
  rom[26918] = 16'hf708;
  rom[26919] = 16'hff29;
  rom[26920] = 16'hff09;
  rom[26921] = 16'hff29;
  rom[26922] = 16'hf708;
  rom[26923] = 16'hff29;
  rom[26924] = 16'hff0a;
  rom[26925] = 16'hff2a;
  rom[26926] = 16'hf70a;
  rom[26927] = 16'hac67;
  rom[26928] = 16'h9a02;
  rom[26929] = 16'hda46;
  rom[26930] = 16'he247;
  rom[26931] = 16'hf1e7;
  rom[26932] = 16'hea27;
  rom[26933] = 16'hda65;
  rom[26934] = 16'hea26;
  rom[26935] = 16'hf227;
  rom[26936] = 16'he1c5;
  rom[26937] = 16'hea27;
  rom[26938] = 16'he207;
  rom[26939] = 16'he228;
  rom[26940] = 16'hda88;
  rom[26941] = 16'haa05;
  rom[26942] = 16'h6960;
  rom[26943] = 16'hc50a;
  rom[26944] = 16'hf6ed;
  rom[26945] = 16'hff0a;
  rom[26946] = 16'hff29;
  rom[26947] = 16'hf72a;
  rom[26948] = 16'hf729;
  rom[26949] = 16'hff49;
  rom[26950] = 16'hef07;
  rom[26951] = 16'hff48;
  rom[26952] = 16'hff28;
  rom[26953] = 16'hff28;
  rom[26954] = 16'hf708;
  rom[26955] = 16'hff29;
  rom[26956] = 16'hff08;
  rom[26957] = 16'hff29;
  rom[26958] = 16'hff08;
  rom[26959] = 16'hff28;
  rom[26960] = 16'hf728;
  rom[26961] = 16'hff08;
  rom[26962] = 16'hf6e9;
  rom[26963] = 16'hf72a;
  rom[26964] = 16'hf72d;
  rom[26965] = 16'hcd2a;
  rom[26966] = 16'h89a1;
  rom[26967] = 16'hca67;
  rom[26968] = 16'hda27;
  rom[26969] = 16'hf247;
  rom[26970] = 16'he226;
  rom[26971] = 16'hea47;
  rom[26972] = 16'hda07;
  rom[26973] = 16'hcb8d;
  rom[26974] = 16'hff5c;
  rom[26975] = 16'hffff;
  rom[26976] = 16'hffff;
  rom[26977] = 16'hffff;
  rom[26978] = 16'hffff;
  rom[26979] = 16'hffff;
  rom[26980] = 16'hffff;
  rom[26981] = 16'hffff;
  rom[26982] = 16'hffff;
  rom[26983] = 16'hffff;
  rom[26984] = 16'hffff;
  rom[26985] = 16'hffff;
  rom[26986] = 16'hffff;
  rom[26987] = 16'hffff;
  rom[26988] = 16'hffff;
  rom[26989] = 16'hffff;
  rom[26990] = 16'hffff;
  rom[26991] = 16'hffff;
  rom[26992] = 16'hffff;
  rom[26993] = 16'hffff;
  rom[26994] = 16'hffff;
  rom[26995] = 16'hffff;
  rom[26996] = 16'hffff;
  rom[26997] = 16'hffff;
  rom[26998] = 16'hffff;
  rom[26999] = 16'hffff;
  rom[27000] = 16'hffff;
  rom[27001] = 16'hffff;
  rom[27002] = 16'hffff;
  rom[27003] = 16'hffff;
  rom[27004] = 16'hffff;
  rom[27005] = 16'hffff;
  rom[27006] = 16'hffff;
  rom[27007] = 16'hffff;
  rom[27008] = 16'hffff;
  rom[27009] = 16'hffbd;
  rom[27010] = 16'hdb6c;
  rom[27011] = 16'hda48;
  rom[27012] = 16'hea07;
  rom[27013] = 16'hea07;
  rom[27014] = 16'hea26;
  rom[27015] = 16'hea26;
  rom[27016] = 16'hf227;
  rom[27017] = 16'hf207;
  rom[27018] = 16'hf227;
  rom[27019] = 16'hf206;
  rom[27020] = 16'hfa07;
  rom[27021] = 16'hf207;
  rom[27022] = 16'hf207;
  rom[27023] = 16'hf207;
  rom[27024] = 16'hf228;
  rom[27025] = 16'hf207;
  rom[27026] = 16'hea27;
  rom[27027] = 16'hea07;
  rom[27028] = 16'hea27;
  rom[27029] = 16'hea26;
  rom[27030] = 16'hea47;
  rom[27031] = 16'hea26;
  rom[27032] = 16'hf227;
  rom[27033] = 16'hf206;
  rom[27034] = 16'hf9e6;
  rom[27035] = 16'hf206;
  rom[27036] = 16'hf227;
  rom[27037] = 16'hf206;
  rom[27038] = 16'hea26;
  rom[27039] = 16'hea06;
  rom[27040] = 16'hf228;
  rom[27041] = 16'hf206;
  rom[27042] = 16'hf227;
  rom[27043] = 16'hea26;
  rom[27044] = 16'hea47;
  rom[27045] = 16'hea26;
  rom[27046] = 16'hea27;
  rom[27047] = 16'hea27;
  rom[27048] = 16'hea28;
  rom[27049] = 16'hea27;
  rom[27050] = 16'hea27;
  rom[27051] = 16'hea07;
  rom[27052] = 16'hf227;
  rom[27053] = 16'hf206;
  rom[27054] = 16'hf226;
  rom[27055] = 16'hea06;
  rom[27056] = 16'hf227;
  rom[27057] = 16'hf206;
  rom[27058] = 16'hf227;
  rom[27059] = 16'hea07;
  rom[27060] = 16'hf227;
  rom[27061] = 16'hea25;
  rom[27062] = 16'hf245;
  rom[27063] = 16'hea25;
  rom[27064] = 16'he267;
  rom[27065] = 16'haa25;
  rom[27066] = 16'h8ac1;
  rom[27067] = 16'hf70c;
  rom[27068] = 16'hf72b;
  rom[27069] = 16'hf709;
  rom[27070] = 16'hff4a;
  rom[27071] = 16'hff29;
  rom[27072] = 16'hff29;
  rom[27073] = 16'hff09;
  rom[27074] = 16'hff0a;
  rom[27075] = 16'hff29;
  rom[27076] = 16'hff29;
  rom[27077] = 16'hff28;
  rom[27078] = 16'hff49;
  rom[27079] = 16'hff4a;
  rom[27080] = 16'hf709;
  rom[27081] = 16'hff49;
  rom[27082] = 16'hf729;
  rom[27083] = 16'hef8b;
  rom[27084] = 16'hee8c;
  rom[27085] = 16'h9ae3;
  rom[27086] = 16'ha204;
  rom[27087] = 16'hc266;
  rom[27088] = 16'hd2a6;
  rom[27089] = 16'hcb23;
  rom[27090] = 16'hfda8;
  rom[27091] = 16'hfec9;
  rom[27092] = 16'hff49;
  rom[27093] = 16'hfea8;
  rom[27094] = 16'hfd86;
  rom[27095] = 16'hcba1;
  rom[27096] = 16'hec44;
  rom[27097] = 16'he423;
  rom[27098] = 16'hdc64;
  rom[27099] = 16'hf5e7;
  rom[27100] = 16'hff28;
  rom[27101] = 16'hff27;
  rom[27102] = 16'hfeca;
  rom[27103] = 16'he464;
  rom[27104] = 16'hdb04;
  rom[27105] = 16'hd265;
  rom[27106] = 16'hd286;
  rom[27107] = 16'h99a2;
  rom[27108] = 16'hab65;
  rom[27109] = 16'hfecc;
  rom[27110] = 16'hfeea;
  rom[27111] = 16'hff49;
  rom[27112] = 16'hf708;
  rom[27113] = 16'hff29;
  rom[27114] = 16'hff2a;
  rom[27115] = 16'hff29;
  rom[27116] = 16'hff29;
  rom[27117] = 16'hff29;
  rom[27118] = 16'hff29;
  rom[27119] = 16'hff08;
  rom[27120] = 16'hff2a;
  rom[27121] = 16'hff28;
  rom[27122] = 16'hff49;
  rom[27123] = 16'hf728;
  rom[27124] = 16'hff29;
  rom[27125] = 16'hf709;
  rom[27126] = 16'hf70c;
  rom[27127] = 16'h8b84;
  rom[27128] = 16'haa24;
  rom[27129] = 16'hda06;
  rom[27130] = 16'hf247;
  rom[27131] = 16'hf207;
  rom[27132] = 16'hf247;
  rom[27133] = 16'he245;
  rom[27134] = 16'hea47;
  rom[27135] = 16'hea07;
  rom[27136] = 16'hf207;
  rom[27137] = 16'hea07;
  rom[27138] = 16'hf227;
  rom[27139] = 16'hea27;
  rom[27140] = 16'hea27;
  rom[27141] = 16'hda87;
  rom[27142] = 16'ha205;
  rom[27143] = 16'h6181;
  rom[27144] = 16'hcd8b;
  rom[27145] = 16'hff2d;
  rom[27146] = 16'hff2a;
  rom[27147] = 16'hf708;
  rom[27148] = 16'hff2a;
  rom[27149] = 16'hf708;
  rom[27150] = 16'hff28;
  rom[27151] = 16'hff28;
  rom[27152] = 16'hff49;
  rom[27153] = 16'hf728;
  rom[27154] = 16'hf729;
  rom[27155] = 16'hff28;
  rom[27156] = 16'hff29;
  rom[27157] = 16'hff29;
  rom[27158] = 16'hf749;
  rom[27159] = 16'hff27;
  rom[27160] = 16'hff08;
  rom[27161] = 16'hff29;
  rom[27162] = 16'hff0a;
  rom[27163] = 16'hf6e9;
  rom[27164] = 16'hff2d;
  rom[27165] = 16'he5cb;
  rom[27166] = 16'h89e2;
  rom[27167] = 16'hba25;
  rom[27168] = 16'hda67;
  rom[27169] = 16'hda25;
  rom[27170] = 16'hea67;
  rom[27171] = 16'he206;
  rom[27172] = 16'hda68;
  rom[27173] = 16'hecd2;
  rom[27174] = 16'hff9e;
  rom[27175] = 16'hffff;
  rom[27176] = 16'hffff;
  rom[27177] = 16'hffff;
  rom[27178] = 16'hffff;
  rom[27179] = 16'hffbf;
  rom[27180] = 16'hffff;
  rom[27181] = 16'hffff;
  rom[27182] = 16'hffff;
  rom[27183] = 16'hffff;
  rom[27184] = 16'hffff;
  rom[27185] = 16'hffff;
  rom[27186] = 16'hffff;
  rom[27187] = 16'hffff;
  rom[27188] = 16'hffff;
  rom[27189] = 16'hffff;
  rom[27190] = 16'hffff;
  rom[27191] = 16'hffff;
  rom[27192] = 16'hffff;
  rom[27193] = 16'hffff;
  rom[27194] = 16'hffff;
  rom[27195] = 16'hffff;
  rom[27196] = 16'hffff;
  rom[27197] = 16'hffff;
  rom[27198] = 16'hffff;
  rom[27199] = 16'hffff;
  rom[27200] = 16'hffff;
  rom[27201] = 16'hffff;
  rom[27202] = 16'hffff;
  rom[27203] = 16'hffff;
  rom[27204] = 16'hffff;
  rom[27205] = 16'hffff;
  rom[27206] = 16'hffff;
  rom[27207] = 16'hffff;
  rom[27208] = 16'hffff;
  rom[27209] = 16'hffdd;
  rom[27210] = 16'hdbee;
  rom[27211] = 16'he269;
  rom[27212] = 16'he207;
  rom[27213] = 16'hf206;
  rom[27214] = 16'hea46;
  rom[27215] = 16'hea46;
  rom[27216] = 16'he206;
  rom[27217] = 16'hf207;
  rom[27218] = 16'hea07;
  rom[27219] = 16'hea26;
  rom[27220] = 16'he206;
  rom[27221] = 16'hf207;
  rom[27222] = 16'hf207;
  rom[27223] = 16'hf207;
  rom[27224] = 16'hea07;
  rom[27225] = 16'hf207;
  rom[27226] = 16'hf207;
  rom[27227] = 16'hf206;
  rom[27228] = 16'hea06;
  rom[27229] = 16'hf226;
  rom[27230] = 16'hea26;
  rom[27231] = 16'hea26;
  rom[27232] = 16'he226;
  rom[27233] = 16'hf226;
  rom[27234] = 16'hea06;
  rom[27235] = 16'hf206;
  rom[27236] = 16'hea06;
  rom[27237] = 16'hf206;
  rom[27238] = 16'hea06;
  rom[27239] = 16'hf207;
  rom[27240] = 16'hea07;
  rom[27241] = 16'hf207;
  rom[27242] = 16'hf206;
  rom[27243] = 16'hea26;
  rom[27244] = 16'hea26;
  rom[27245] = 16'hea07;
  rom[27246] = 16'hea07;
  rom[27247] = 16'hea27;
  rom[27248] = 16'hea27;
  rom[27249] = 16'hea27;
  rom[27250] = 16'hea27;
  rom[27251] = 16'hf207;
  rom[27252] = 16'hea06;
  rom[27253] = 16'hf206;
  rom[27254] = 16'hf206;
  rom[27255] = 16'hf206;
  rom[27256] = 16'he226;
  rom[27257] = 16'hea26;
  rom[27258] = 16'hea06;
  rom[27259] = 16'hf208;
  rom[27260] = 16'hea06;
  rom[27261] = 16'hea26;
  rom[27262] = 16'hf225;
  rom[27263] = 16'hf226;
  rom[27264] = 16'he247;
  rom[27265] = 16'hb225;
  rom[27266] = 16'h7a00;
  rom[27267] = 16'hff0e;
  rom[27268] = 16'hf70b;
  rom[27269] = 16'hf729;
  rom[27270] = 16'hf708;
  rom[27271] = 16'hff29;
  rom[27272] = 16'hf709;
  rom[27273] = 16'hff09;
  rom[27274] = 16'hff09;
  rom[27275] = 16'hff29;
  rom[27276] = 16'hf707;
  rom[27277] = 16'hff48;
  rom[27278] = 16'hf708;
  rom[27279] = 16'hf729;
  rom[27280] = 16'hf709;
  rom[27281] = 16'hff2a;
  rom[27282] = 16'hf6e9;
  rom[27283] = 16'hf74c;
  rom[27284] = 16'hbce6;
  rom[27285] = 16'h89c1;
  rom[27286] = 16'hca87;
  rom[27287] = 16'hda88;
  rom[27288] = 16'hd284;
  rom[27289] = 16'hdc25;
  rom[27290] = 16'hfe29;
  rom[27291] = 16'hfec9;
  rom[27292] = 16'hfe47;
  rom[27293] = 16'hfd26;
  rom[27294] = 16'hd322;
  rom[27295] = 16'hd2e3;
  rom[27296] = 16'hec06;
  rom[27297] = 16'he3e5;
  rom[27298] = 16'hc322;
  rom[27299] = 16'hcb82;
  rom[27300] = 16'hfd66;
  rom[27301] = 16'hfe69;
  rom[27302] = 16'hfea9;
  rom[27303] = 16'hfe2a;
  rom[27304] = 16'hd363;
  rom[27305] = 16'hda84;
  rom[27306] = 16'hd246;
  rom[27307] = 16'hca86;
  rom[27308] = 16'h9201;
  rom[27309] = 16'hd569;
  rom[27310] = 16'hf70c;
  rom[27311] = 16'hf6e9;
  rom[27312] = 16'hff6a;
  rom[27313] = 16'hff4a;
  rom[27314] = 16'hf6e9;
  rom[27315] = 16'hff2a;
  rom[27316] = 16'hf72a;
  rom[27317] = 16'hff29;
  rom[27318] = 16'hf709;
  rom[27319] = 16'hff4a;
  rom[27320] = 16'hf709;
  rom[27321] = 16'hff4a;
  rom[27322] = 16'hf708;
  rom[27323] = 16'hf728;
  rom[27324] = 16'hf708;
  rom[27325] = 16'hff2a;
  rom[27326] = 16'hf6ec;
  rom[27327] = 16'h7ae2;
  rom[27328] = 16'ha9e4;
  rom[27329] = 16'hea27;
  rom[27330] = 16'hea07;
  rom[27331] = 16'hf207;
  rom[27332] = 16'hea05;
  rom[27333] = 16'hea45;
  rom[27334] = 16'hea26;
  rom[27335] = 16'hf227;
  rom[27336] = 16'he9e7;
  rom[27337] = 16'hf207;
  rom[27338] = 16'hea27;
  rom[27339] = 16'hf227;
  rom[27340] = 16'hea05;
  rom[27341] = 16'he226;
  rom[27342] = 16'hcaa8;
  rom[27343] = 16'h6941;
  rom[27344] = 16'h7b04;
  rom[27345] = 16'hf6ee;
  rom[27346] = 16'hf70a;
  rom[27347] = 16'hff29;
  rom[27348] = 16'hff28;
  rom[27349] = 16'hff49;
  rom[27350] = 16'hff29;
  rom[27351] = 16'hf708;
  rom[27352] = 16'hf728;
  rom[27353] = 16'hf748;
  rom[27354] = 16'hf728;
  rom[27355] = 16'hff49;
  rom[27356] = 16'hf708;
  rom[27357] = 16'hff29;
  rom[27358] = 16'hf728;
  rom[27359] = 16'hff28;
  rom[27360] = 16'hf6e8;
  rom[27361] = 16'hff0a;
  rom[27362] = 16'hfeea;
  rom[27363] = 16'hff0a;
  rom[27364] = 16'hf70b;
  rom[27365] = 16'hee2c;
  rom[27366] = 16'h8a42;
  rom[27367] = 16'haa25;
  rom[27368] = 16'hd246;
  rom[27369] = 16'hda45;
  rom[27370] = 16'he225;
  rom[27371] = 16'he247;
  rom[27372] = 16'hd2ca;
  rom[27373] = 16'hfdf7;
  rom[27374] = 16'hff9e;
  rom[27375] = 16'hffff;
  rom[27376] = 16'hfffe;
  rom[27377] = 16'hffff;
  rom[27378] = 16'hffff;
  rom[27379] = 16'hffdf;
  rom[27380] = 16'hffdf;
  rom[27381] = 16'hffff;
  rom[27382] = 16'hffff;
  rom[27383] = 16'hffff;
  rom[27384] = 16'hffff;
  rom[27385] = 16'hffff;
  rom[27386] = 16'hffff;
  rom[27387] = 16'hffff;
  rom[27388] = 16'hffff;
  rom[27389] = 16'hffff;
  rom[27390] = 16'hffff;
  rom[27391] = 16'hffff;
  rom[27392] = 16'hffff;
  rom[27393] = 16'hffff;
  rom[27394] = 16'hffff;
  rom[27395] = 16'hffff;
  rom[27396] = 16'hffff;
  rom[27397] = 16'hffff;
  rom[27398] = 16'hffff;
  rom[27399] = 16'hffff;
  rom[27400] = 16'hffff;
  rom[27401] = 16'hffff;
  rom[27402] = 16'hffff;
  rom[27403] = 16'hffff;
  rom[27404] = 16'hffff;
  rom[27405] = 16'hffff;
  rom[27406] = 16'hffff;
  rom[27407] = 16'hffff;
  rom[27408] = 16'hffff;
  rom[27409] = 16'hffbd;
  rom[27410] = 16'hf4b1;
  rom[27411] = 16'hda89;
  rom[27412] = 16'he9e6;
  rom[27413] = 16'hf226;
  rom[27414] = 16'hea47;
  rom[27415] = 16'he246;
  rom[27416] = 16'hea27;
  rom[27417] = 16'hf207;
  rom[27418] = 16'hf227;
  rom[27419] = 16'hea26;
  rom[27420] = 16'hea46;
  rom[27421] = 16'hea07;
  rom[27422] = 16'hf228;
  rom[27423] = 16'hf207;
  rom[27424] = 16'hf227;
  rom[27425] = 16'hf207;
  rom[27426] = 16'hf228;
  rom[27427] = 16'hf206;
  rom[27428] = 16'hf226;
  rom[27429] = 16'hf206;
  rom[27430] = 16'hea47;
  rom[27431] = 16'hea26;
  rom[27432] = 16'hea46;
  rom[27433] = 16'hea26;
  rom[27434] = 16'hea47;
  rom[27435] = 16'hea26;
  rom[27436] = 16'hea46;
  rom[27437] = 16'hea26;
  rom[27438] = 16'hea28;
  rom[27439] = 16'hea07;
  rom[27440] = 16'hf228;
  rom[27441] = 16'hf208;
  rom[27442] = 16'hf208;
  rom[27443] = 16'hf208;
  rom[27444] = 16'hf228;
  rom[27445] = 16'hf206;
  rom[27446] = 16'hf227;
  rom[27447] = 16'hf206;
  rom[27448] = 16'hf226;
  rom[27449] = 16'hf206;
  rom[27450] = 16'hf227;
  rom[27451] = 16'hf206;
  rom[27452] = 16'hf226;
  rom[27453] = 16'hf206;
  rom[27454] = 16'hf227;
  rom[27455] = 16'hea26;
  rom[27456] = 16'hea46;
  rom[27457] = 16'he246;
  rom[27458] = 16'hea47;
  rom[27459] = 16'hea07;
  rom[27460] = 16'hea27;
  rom[27461] = 16'hea26;
  rom[27462] = 16'hf246;
  rom[27463] = 16'hf206;
  rom[27464] = 16'hea48;
  rom[27465] = 16'hc246;
  rom[27466] = 16'h81c1;
  rom[27467] = 16'hfece;
  rom[27468] = 16'hff0b;
  rom[27469] = 16'hff09;
  rom[27470] = 16'hff29;
  rom[27471] = 16'hff28;
  rom[27472] = 16'hff28;
  rom[27473] = 16'hf728;
  rom[27474] = 16'hff29;
  rom[27475] = 16'hff28;
  rom[27476] = 16'hff48;
  rom[27477] = 16'hf729;
  rom[27478] = 16'hff2a;
  rom[27479] = 16'hef09;
  rom[27480] = 16'hff4b;
  rom[27481] = 16'hff2a;
  rom[27482] = 16'hfeeb;
  rom[27483] = 16'heeac;
  rom[27484] = 16'hab63;
  rom[27485] = 16'haa03;
  rom[27486] = 16'hd206;
  rom[27487] = 16'hda67;
  rom[27488] = 16'hd2a4;
  rom[27489] = 16'hfd69;
  rom[27490] = 16'hfe6b;
  rom[27491] = 16'hfdc9;
  rom[27492] = 16'he404;
  rom[27493] = 16'hcaa2;
  rom[27494] = 16'hd2c4;
  rom[27495] = 16'hd325;
  rom[27496] = 16'hfd0b;
  rom[27497] = 16'heca9;
  rom[27498] = 16'hd2e4;
  rom[27499] = 16'hd2a3;
  rom[27500] = 16'hdae3;
  rom[27501] = 16'hec66;
  rom[27502] = 16'hfdc9;
  rom[27503] = 16'hfe6c;
  rom[27504] = 16'hf4e8;
  rom[27505] = 16'hca62;
  rom[27506] = 16'he2a7;
  rom[27507] = 16'hd287;
  rom[27508] = 16'haa43;
  rom[27509] = 16'habc5;
  rom[27510] = 16'hff10;
  rom[27511] = 16'hfecd;
  rom[27512] = 16'hfeed;
  rom[27513] = 16'hf70c;
  rom[27514] = 16'hff2c;
  rom[27515] = 16'hff2c;
  rom[27516] = 16'hff0c;
  rom[27517] = 16'hf70b;
  rom[27518] = 16'hff2b;
  rom[27519] = 16'hf70b;
  rom[27520] = 16'hff4b;
  rom[27521] = 16'hf70a;
  rom[27522] = 16'hf70a;
  rom[27523] = 16'hf72a;
  rom[27524] = 16'hf72b;
  rom[27525] = 16'hf72c;
  rom[27526] = 16'hff0f;
  rom[27527] = 16'h7a62;
  rom[27528] = 16'hba26;
  rom[27529] = 16'hea07;
  rom[27530] = 16'hf208;
  rom[27531] = 16'hea07;
  rom[27532] = 16'hea26;
  rom[27533] = 16'hea26;
  rom[27534] = 16'hea27;
  rom[27535] = 16'hf207;
  rom[27536] = 16'hf227;
  rom[27537] = 16'hf206;
  rom[27538] = 16'hea27;
  rom[27539] = 16'hf206;
  rom[27540] = 16'hf226;
  rom[27541] = 16'hea05;
  rom[27542] = 16'hd2a8;
  rom[27543] = 16'h9aa6;
  rom[27544] = 16'h7263;
  rom[27545] = 16'he6ac;
  rom[27546] = 16'hf70a;
  rom[27547] = 16'hff48;
  rom[27548] = 16'hff49;
  rom[27549] = 16'hff29;
  rom[27550] = 16'hff2a;
  rom[27551] = 16'hff2a;
  rom[27552] = 16'hff2a;
  rom[27553] = 16'hf709;
  rom[27554] = 16'hf72a;
  rom[27555] = 16'hff29;
  rom[27556] = 16'hff2a;
  rom[27557] = 16'hff29;
  rom[27558] = 16'hff29;
  rom[27559] = 16'hff28;
  rom[27560] = 16'hff09;
  rom[27561] = 16'hfee9;
  rom[27562] = 16'hff2a;
  rom[27563] = 16'hff09;
  rom[27564] = 16'hff6b;
  rom[27565] = 16'hee6c;
  rom[27566] = 16'h92a3;
  rom[27567] = 16'ha204;
  rom[27568] = 16'hda88;
  rom[27569] = 16'he226;
  rom[27570] = 16'hea27;
  rom[27571] = 16'hd247;
  rom[27572] = 16'hd38d;
  rom[27573] = 16'hfeda;
  rom[27574] = 16'hffff;
  rom[27575] = 16'hffff;
  rom[27576] = 16'hffff;
  rom[27577] = 16'hffff;
  rom[27578] = 16'hffff;
  rom[27579] = 16'hffff;
  rom[27580] = 16'hffff;
  rom[27581] = 16'hffff;
  rom[27582] = 16'hffff;
  rom[27583] = 16'hffff;
  rom[27584] = 16'hffff;
  rom[27585] = 16'hffff;
  rom[27586] = 16'hffff;
  rom[27587] = 16'hffff;
  rom[27588] = 16'hffff;
  rom[27589] = 16'hffff;
  rom[27590] = 16'hffff;
  rom[27591] = 16'hffff;
  rom[27592] = 16'hffff;
  rom[27593] = 16'hffff;
  rom[27594] = 16'hffff;
  rom[27595] = 16'hffff;
  rom[27596] = 16'hffff;
  rom[27597] = 16'hffff;
  rom[27598] = 16'hffff;
  rom[27599] = 16'hffff;
  rom[27600] = 16'hffff;
  rom[27601] = 16'hffff;
  rom[27602] = 16'hffff;
  rom[27603] = 16'hffff;
  rom[27604] = 16'hffff;
  rom[27605] = 16'hffff;
  rom[27606] = 16'hffff;
  rom[27607] = 16'hffdf;
  rom[27608] = 16'hffff;
  rom[27609] = 16'hffde;
  rom[27610] = 16'hf553;
  rom[27611] = 16'hdaa9;
  rom[27612] = 16'he1e6;
  rom[27613] = 16'hf226;
  rom[27614] = 16'hea25;
  rom[27615] = 16'hea46;
  rom[27616] = 16'hea27;
  rom[27617] = 16'hea07;
  rom[27618] = 16'he206;
  rom[27619] = 16'hea26;
  rom[27620] = 16'hea26;
  rom[27621] = 16'hea27;
  rom[27622] = 16'hea07;
  rom[27623] = 16'hf207;
  rom[27624] = 16'hf207;
  rom[27625] = 16'hf207;
  rom[27626] = 16'hea07;
  rom[27627] = 16'hf206;
  rom[27628] = 16'hf206;
  rom[27629] = 16'hf226;
  rom[27630] = 16'he226;
  rom[27631] = 16'hea26;
  rom[27632] = 16'hea26;
  rom[27633] = 16'hea26;
  rom[27634] = 16'he227;
  rom[27635] = 16'hea27;
  rom[27636] = 16'hea27;
  rom[27637] = 16'hea27;
  rom[27638] = 16'he207;
  rom[27639] = 16'hea07;
  rom[27640] = 16'hf207;
  rom[27641] = 16'hf208;
  rom[27642] = 16'hea08;
  rom[27643] = 16'hf208;
  rom[27644] = 16'hf207;
  rom[27645] = 16'hf206;
  rom[27646] = 16'hea26;
  rom[27647] = 16'hf206;
  rom[27648] = 16'hf206;
  rom[27649] = 16'hf206;
  rom[27650] = 16'hea06;
  rom[27651] = 16'hf206;
  rom[27652] = 16'hf206;
  rom[27653] = 16'hf207;
  rom[27654] = 16'hea07;
  rom[27655] = 16'hea27;
  rom[27656] = 16'he226;
  rom[27657] = 16'he246;
  rom[27658] = 16'he226;
  rom[27659] = 16'hea27;
  rom[27660] = 16'hea27;
  rom[27661] = 16'hea26;
  rom[27662] = 16'hea45;
  rom[27663] = 16'hf206;
  rom[27664] = 16'hea08;
  rom[27665] = 16'hca46;
  rom[27666] = 16'h7941;
  rom[27667] = 16'he5ec;
  rom[27668] = 16'hf70b;
  rom[27669] = 16'hff29;
  rom[27670] = 16'hf728;
  rom[27671] = 16'hf707;
  rom[27672] = 16'hf728;
  rom[27673] = 16'hff6a;
  rom[27674] = 16'hf749;
  rom[27675] = 16'heee8;
  rom[27676] = 16'hf70a;
  rom[27677] = 16'hff0b;
  rom[27678] = 16'hff2c;
  rom[27679] = 16'hff4c;
  rom[27680] = 16'he68a;
  rom[27681] = 16'hff0d;
  rom[27682] = 16'hf6ce;
  rom[27683] = 16'hd54b;
  rom[27684] = 16'h89e1;
  rom[27685] = 16'hca46;
  rom[27686] = 16'heaa8;
  rom[27687] = 16'hda45;
  rom[27688] = 16'hfc49;
  rom[27689] = 16'hfdeb;
  rom[27690] = 16'hfd27;
  rom[27691] = 16'hd322;
  rom[27692] = 16'hdaa2;
  rom[27693] = 16'he264;
  rom[27694] = 16'hd284;
  rom[27695] = 16'hec08;
  rom[27696] = 16'hfe2d;
  rom[27697] = 16'hfe0d;
  rom[27698] = 16'hebe7;
  rom[27699] = 16'he284;
  rom[27700] = 16'he265;
  rom[27701] = 16'hd262;
  rom[27702] = 16'hdbc3;
  rom[27703] = 16'hfdca;
  rom[27704] = 16'hfdeb;
  rom[27705] = 16'he3a6;
  rom[27706] = 16'hca65;
  rom[27707] = 16'hda47;
  rom[27708] = 16'ha1c3;
  rom[27709] = 16'h8a43;
  rom[27710] = 16'hd4ea;
  rom[27711] = 16'hed8e;
  rom[27712] = 16'hdd2b;
  rom[27713] = 16'hd56a;
  rom[27714] = 16'hd56a;
  rom[27715] = 16'hd56a;
  rom[27716] = 16'hdd8a;
  rom[27717] = 16'hddcb;
  rom[27718] = 16'he60b;
  rom[27719] = 16'hee2b;
  rom[27720] = 16'hddea;
  rom[27721] = 16'hf6ac;
  rom[27722] = 16'hff4e;
  rom[27723] = 16'hff2e;
  rom[27724] = 16'hf6cd;
  rom[27725] = 16'hf6ce;
  rom[27726] = 16'hcd6b;
  rom[27727] = 16'h71a1;
  rom[27728] = 16'hb9e6;
  rom[27729] = 16'hf228;
  rom[27730] = 16'he9e7;
  rom[27731] = 16'hea27;
  rom[27732] = 16'hea26;
  rom[27733] = 16'hea26;
  rom[27734] = 16'he206;
  rom[27735] = 16'hea07;
  rom[27736] = 16'hea07;
  rom[27737] = 16'hea26;
  rom[27738] = 16'hea06;
  rom[27739] = 16'hf206;
  rom[27740] = 16'hf206;
  rom[27741] = 16'hea26;
  rom[27742] = 16'hd287;
  rom[27743] = 16'h8a03;
  rom[27744] = 16'h8b46;
  rom[27745] = 16'hff0e;
  rom[27746] = 16'hff6b;
  rom[27747] = 16'hff68;
  rom[27748] = 16'hf727;
  rom[27749] = 16'hf708;
  rom[27750] = 16'heec8;
  rom[27751] = 16'hff2a;
  rom[27752] = 16'hff2a;
  rom[27753] = 16'hff2a;
  rom[27754] = 16'hf70a;
  rom[27755] = 16'hff29;
  rom[27756] = 16'hf709;
  rom[27757] = 16'hff29;
  rom[27758] = 16'hf708;
  rom[27759] = 16'hff48;
  rom[27760] = 16'hff08;
  rom[27761] = 16'hff29;
  rom[27762] = 16'hf709;
  rom[27763] = 16'hf728;
  rom[27764] = 16'hf72a;
  rom[27765] = 16'he68c;
  rom[27766] = 16'h8ac2;
  rom[27767] = 16'h9a05;
  rom[27768] = 16'hd227;
  rom[27769] = 16'hf207;
  rom[27770] = 16'he206;
  rom[27771] = 16'hca89;
  rom[27772] = 16'hf594;
  rom[27773] = 16'hff7c;
  rom[27774] = 16'hf7fe;
  rom[27775] = 16'hffff;
  rom[27776] = 16'hffff;
  rom[27777] = 16'hffff;
  rom[27778] = 16'hffff;
  rom[27779] = 16'hffff;
  rom[27780] = 16'hffff;
  rom[27781] = 16'hffff;
  rom[27782] = 16'hffff;
  rom[27783] = 16'hffff;
  rom[27784] = 16'hffff;
  rom[27785] = 16'hffff;
  rom[27786] = 16'hffff;
  rom[27787] = 16'hffff;
  rom[27788] = 16'hffff;
  rom[27789] = 16'hffff;
  rom[27790] = 16'hffff;
  rom[27791] = 16'hffff;
  rom[27792] = 16'hffff;
  rom[27793] = 16'hffff;
  rom[27794] = 16'hffff;
  rom[27795] = 16'hffff;
  rom[27796] = 16'hffff;
  rom[27797] = 16'hffff;
  rom[27798] = 16'hffff;
  rom[27799] = 16'hffff;
  rom[27800] = 16'hffff;
  rom[27801] = 16'hffff;
  rom[27802] = 16'hffff;
  rom[27803] = 16'hffff;
  rom[27804] = 16'hffff;
  rom[27805] = 16'hffff;
  rom[27806] = 16'hffff;
  rom[27807] = 16'hffff;
  rom[27808] = 16'hffff;
  rom[27809] = 16'hfffe;
  rom[27810] = 16'hfe57;
  rom[27811] = 16'hd30b;
  rom[27812] = 16'he228;
  rom[27813] = 16'hf227;
  rom[27814] = 16'hea26;
  rom[27815] = 16'hea46;
  rom[27816] = 16'hea47;
  rom[27817] = 16'hea07;
  rom[27818] = 16'hea27;
  rom[27819] = 16'hea26;
  rom[27820] = 16'hea47;
  rom[27821] = 16'hea27;
  rom[27822] = 16'hea27;
  rom[27823] = 16'hf207;
  rom[27824] = 16'hf228;
  rom[27825] = 16'hf207;
  rom[27826] = 16'hf227;
  rom[27827] = 16'hea06;
  rom[27828] = 16'hf227;
  rom[27829] = 16'hea06;
  rom[27830] = 16'hea46;
  rom[27831] = 16'hea26;
  rom[27832] = 16'hea47;
  rom[27833] = 16'hea26;
  rom[27834] = 16'hea27;
  rom[27835] = 16'hea27;
  rom[27836] = 16'hf228;
  rom[27837] = 16'hea07;
  rom[27838] = 16'hf227;
  rom[27839] = 16'hf207;
  rom[27840] = 16'hf227;
  rom[27841] = 16'hf207;
  rom[27842] = 16'hf227;
  rom[27843] = 16'hea27;
  rom[27844] = 16'hf227;
  rom[27845] = 16'hea26;
  rom[27846] = 16'hea46;
  rom[27847] = 16'hea26;
  rom[27848] = 16'hf227;
  rom[27849] = 16'hea26;
  rom[27850] = 16'hf226;
  rom[27851] = 16'hea26;
  rom[27852] = 16'hf227;
  rom[27853] = 16'hf206;
  rom[27854] = 16'hf227;
  rom[27855] = 16'hea07;
  rom[27856] = 16'hf227;
  rom[27857] = 16'hea46;
  rom[27858] = 16'hea27;
  rom[27859] = 16'hea27;
  rom[27860] = 16'hea27;
  rom[27861] = 16'hea26;
  rom[27862] = 16'hf245;
  rom[27863] = 16'hea06;
  rom[27864] = 16'hea49;
  rom[27865] = 16'hca68;
  rom[27866] = 16'h8162;
  rom[27867] = 16'hbca8;
  rom[27868] = 16'hff0d;
  rom[27869] = 16'heeea;
  rom[27870] = 16'hff2a;
  rom[27871] = 16'hf72a;
  rom[27872] = 16'hff2b;
  rom[27873] = 16'hf70c;
  rom[27874] = 16'hf70d;
  rom[27875] = 16'hf6cc;
  rom[27876] = 16'hf66c;
  rom[27877] = 16'hf60c;
  rom[27878] = 16'he58b;
  rom[27879] = 16'hc4c7;
  rom[27880] = 16'hbc87;
  rom[27881] = 16'hb428;
  rom[27882] = 16'ha387;
  rom[27883] = 16'h8243;
  rom[27884] = 16'h9142;
  rom[27885] = 16'hd226;
  rom[27886] = 16'he247;
  rom[27887] = 16'heb07;
  rom[27888] = 16'hfd0b;
  rom[27889] = 16'hecc7;
  rom[27890] = 16'hd3a2;
  rom[27891] = 16'hcae1;
  rom[27892] = 16'he2a4;
  rom[27893] = 16'hda44;
  rom[27894] = 16'heb46;
  rom[27895] = 16'hfdaa;
  rom[27896] = 16'hff0b;
  rom[27897] = 16'hfeca;
  rom[27898] = 16'hfd28;
  rom[27899] = 16'he2e4;
  rom[27900] = 16'hea66;
  rom[27901] = 16'hda63;
  rom[27902] = 16'hdb02;
  rom[27903] = 16'hcb42;
  rom[27904] = 16'hfd09;
  rom[27905] = 16'hfcca;
  rom[27906] = 16'hdae7;
  rom[27907] = 16'he268;
  rom[27908] = 16'hca69;
  rom[27909] = 16'h7101;
  rom[27910] = 16'h7962;
  rom[27911] = 16'h81a3;
  rom[27912] = 16'h89c4;
  rom[27913] = 16'h81a2;
  rom[27914] = 16'h89e2;
  rom[27915] = 16'h81c1;
  rom[27916] = 16'h81c2;
  rom[27917] = 16'h81e1;
  rom[27918] = 16'h89e1;
  rom[27919] = 16'h8201;
  rom[27920] = 16'h9aa3;
  rom[27921] = 16'h9ae4;
  rom[27922] = 16'hab25;
  rom[27923] = 16'hb3a6;
  rom[27924] = 16'hbc27;
  rom[27925] = 16'hb468;
  rom[27926] = 16'ha3a7;
  rom[27927] = 16'h8182;
  rom[27928] = 16'hd249;
  rom[27929] = 16'hea08;
  rom[27930] = 16'hf227;
  rom[27931] = 16'hea47;
  rom[27932] = 16'hea47;
  rom[27933] = 16'hea26;
  rom[27934] = 16'hf227;
  rom[27935] = 16'hea07;
  rom[27936] = 16'hea27;
  rom[27937] = 16'hea06;
  rom[27938] = 16'hf247;
  rom[27939] = 16'hf206;
  rom[27940] = 16'hf227;
  rom[27941] = 16'hea26;
  rom[27942] = 16'hd267;
  rom[27943] = 16'h8182;
  rom[27944] = 16'hac09;
  rom[27945] = 16'hf6ce;
  rom[27946] = 16'hf70a;
  rom[27947] = 16'hf727;
  rom[27948] = 16'hf748;
  rom[27949] = 16'hff49;
  rom[27950] = 16'hff4a;
  rom[27951] = 16'hff09;
  rom[27952] = 16'hff29;
  rom[27953] = 16'hff09;
  rom[27954] = 16'hff29;
  rom[27955] = 16'hff29;
  rom[27956] = 16'hff29;
  rom[27957] = 16'hff29;
  rom[27958] = 16'hff29;
  rom[27959] = 16'hff28;
  rom[27960] = 16'hff2a;
  rom[27961] = 16'hff29;
  rom[27962] = 16'hff29;
  rom[27963] = 16'hf748;
  rom[27964] = 16'hf74a;
  rom[27965] = 16'hee8c;
  rom[27966] = 16'h9b04;
  rom[27967] = 16'ha1c4;
  rom[27968] = 16'hda69;
  rom[27969] = 16'he1c6;
  rom[27970] = 16'hda49;
  rom[27971] = 16'hdbce;
  rom[27972] = 16'hff1b;
  rom[27973] = 16'hffdd;
  rom[27974] = 16'hffff;
  rom[27975] = 16'hffff;
  rom[27976] = 16'hffff;
  rom[27977] = 16'hffff;
  rom[27978] = 16'hffff;
  rom[27979] = 16'hffff;
  rom[27980] = 16'hffff;
  rom[27981] = 16'hffff;
  rom[27982] = 16'hffff;
  rom[27983] = 16'hffff;
  rom[27984] = 16'hffff;
  rom[27985] = 16'hffff;
  rom[27986] = 16'hffff;
  rom[27987] = 16'hffff;
  rom[27988] = 16'hffff;
  rom[27989] = 16'hffff;
  rom[27990] = 16'hffff;
  rom[27991] = 16'hffff;
  rom[27992] = 16'hffff;
  rom[27993] = 16'hffff;
  rom[27994] = 16'hffff;
  rom[27995] = 16'hffff;
  rom[27996] = 16'hffff;
  rom[27997] = 16'hffff;
  rom[27998] = 16'hffff;
  rom[27999] = 16'hffff;
  rom[28000] = 16'hffff;
  rom[28001] = 16'hffff;
  rom[28002] = 16'hffff;
  rom[28003] = 16'hffff;
  rom[28004] = 16'hffff;
  rom[28005] = 16'hffff;
  rom[28006] = 16'hffff;
  rom[28007] = 16'hffff;
  rom[28008] = 16'hffff;
  rom[28009] = 16'hfffe;
  rom[28010] = 16'hfed9;
  rom[28011] = 16'hd34c;
  rom[28012] = 16'hda27;
  rom[28013] = 16'hf227;
  rom[28014] = 16'hea05;
  rom[28015] = 16'hf226;
  rom[28016] = 16'he226;
  rom[28017] = 16'hf207;
  rom[28018] = 16'hea06;
  rom[28019] = 16'hea26;
  rom[28020] = 16'hea06;
  rom[28021] = 16'hea07;
  rom[28022] = 16'hea07;
  rom[28023] = 16'hf207;
  rom[28024] = 16'hea07;
  rom[28025] = 16'hea07;
  rom[28026] = 16'hea06;
  rom[28027] = 16'hea06;
  rom[28028] = 16'he206;
  rom[28029] = 16'hea26;
  rom[28030] = 16'hea26;
  rom[28031] = 16'hea26;
  rom[28032] = 16'he226;
  rom[28033] = 16'hea26;
  rom[28034] = 16'hea07;
  rom[28035] = 16'hf207;
  rom[28036] = 16'hea07;
  rom[28037] = 16'hf207;
  rom[28038] = 16'hf206;
  rom[28039] = 16'hf206;
  rom[28040] = 16'hea06;
  rom[28041] = 16'hea26;
  rom[28042] = 16'hea26;
  rom[28043] = 16'hea26;
  rom[28044] = 16'he226;
  rom[28045] = 16'hea26;
  rom[28046] = 16'he246;
  rom[28047] = 16'hea26;
  rom[28048] = 16'he226;
  rom[28049] = 16'hea26;
  rom[28050] = 16'hea26;
  rom[28051] = 16'hea26;
  rom[28052] = 16'he226;
  rom[28053] = 16'hea26;
  rom[28054] = 16'hea07;
  rom[28055] = 16'hf207;
  rom[28056] = 16'hea06;
  rom[28057] = 16'hf226;
  rom[28058] = 16'hea06;
  rom[28059] = 16'hf207;
  rom[28060] = 16'hea06;
  rom[28061] = 16'hea26;
  rom[28062] = 16'hea26;
  rom[28063] = 16'hf227;
  rom[28064] = 16'he228;
  rom[28065] = 16'hca88;
  rom[28066] = 16'h7982;
  rom[28067] = 16'h8b65;
  rom[28068] = 16'hf70e;
  rom[28069] = 16'hf70d;
  rom[28070] = 16'hff2c;
  rom[28071] = 16'hfeed;
  rom[28072] = 16'hee4b;
  rom[28073] = 16'hdd8a;
  rom[28074] = 16'hc4c8;
  rom[28075] = 16'hb3e6;
  rom[28076] = 16'h92a2;
  rom[28077] = 16'h81c2;
  rom[28078] = 16'h89a1;
  rom[28079] = 16'h89c1;
  rom[28080] = 16'h8a02;
  rom[28081] = 16'h89e3;
  rom[28082] = 16'h9245;
  rom[28083] = 16'h7963;
  rom[28084] = 16'h9184;
  rom[28085] = 16'hda68;
  rom[28086] = 16'hda67;
  rom[28087] = 16'hfc0a;
  rom[28088] = 16'hfd0b;
  rom[28089] = 16'hec26;
  rom[28090] = 16'he3c4;
  rom[28091] = 16'hdb24;
  rom[28092] = 16'hdaa4;
  rom[28093] = 16'hd284;
  rom[28094] = 16'hec87;
  rom[28095] = 16'hfec9;
  rom[28096] = 16'hff66;
  rom[28097] = 16'hff67;
  rom[28098] = 16'hfe68;
  rom[28099] = 16'hebe5;
  rom[28100] = 16'hd284;
  rom[28101] = 16'he2a5;
  rom[28102] = 16'hdae3;
  rom[28103] = 16'heb85;
  rom[28104] = 16'hfc47;
  rom[28105] = 16'hfd0b;
  rom[28106] = 16'hebca;
  rom[28107] = 16'hd227;
  rom[28108] = 16'hca49;
  rom[28109] = 16'h9165;
  rom[28110] = 16'h9964;
  rom[28111] = 16'hc288;
  rom[28112] = 16'hcaa7;
  rom[28113] = 16'hc267;
  rom[28114] = 16'hc287;
  rom[28115] = 16'hca88;
  rom[28116] = 16'hc267;
  rom[28117] = 16'hca66;
  rom[28118] = 16'hc246;
  rom[28119] = 16'hc266;
  rom[28120] = 16'hc266;
  rom[28121] = 16'hc287;
  rom[28122] = 16'hba45;
  rom[28123] = 16'hb224;
  rom[28124] = 16'h91e2;
  rom[28125] = 16'h8202;
  rom[28126] = 16'h6120;
  rom[28127] = 16'h8122;
  rom[28128] = 16'hda68;
  rom[28129] = 16'he1c7;
  rom[28130] = 16'hf207;
  rom[28131] = 16'hea47;
  rom[28132] = 16'he226;
  rom[28133] = 16'hf226;
  rom[28134] = 16'hf206;
  rom[28135] = 16'hea27;
  rom[28136] = 16'hea27;
  rom[28137] = 16'hf207;
  rom[28138] = 16'hf206;
  rom[28139] = 16'hf206;
  rom[28140] = 16'hea06;
  rom[28141] = 16'hea27;
  rom[28142] = 16'hda87;
  rom[28143] = 16'h7900;
  rom[28144] = 16'hb429;
  rom[28145] = 16'hff10;
  rom[28146] = 16'hef0c;
  rom[28147] = 16'hf729;
  rom[28148] = 16'hef08;
  rom[28149] = 16'hf709;
  rom[28150] = 16'hef07;
  rom[28151] = 16'hff29;
  rom[28152] = 16'hff28;
  rom[28153] = 16'hff48;
  rom[28154] = 16'hff28;
  rom[28155] = 16'hff28;
  rom[28156] = 16'hf708;
  rom[28157] = 16'hff29;
  rom[28158] = 16'hff09;
  rom[28159] = 16'hf729;
  rom[28160] = 16'hf709;
  rom[28161] = 16'hff09;
  rom[28162] = 16'hff08;
  rom[28163] = 16'hf748;
  rom[28164] = 16'hef29;
  rom[28165] = 16'hee4b;
  rom[28166] = 16'h9242;
  rom[28167] = 16'ha9a4;
  rom[28168] = 16'hda89;
  rom[28169] = 16'hd207;
  rom[28170] = 16'hd30b;
  rom[28171] = 16'hfe18;
  rom[28172] = 16'hff9d;
  rom[28173] = 16'hffff;
  rom[28174] = 16'hffff;
  rom[28175] = 16'hffff;
  rom[28176] = 16'hffff;
  rom[28177] = 16'hffff;
  rom[28178] = 16'hffff;
  rom[28179] = 16'hffff;
  rom[28180] = 16'hffff;
  rom[28181] = 16'hffff;
  rom[28182] = 16'hffff;
  rom[28183] = 16'hffff;
  rom[28184] = 16'hffff;
  rom[28185] = 16'hffff;
  rom[28186] = 16'hffff;
  rom[28187] = 16'hffff;
  rom[28188] = 16'hffff;
  rom[28189] = 16'hffff;
  rom[28190] = 16'hffff;
  rom[28191] = 16'hffff;
  rom[28192] = 16'hffff;
  rom[28193] = 16'hffff;
  rom[28194] = 16'hffff;
  rom[28195] = 16'hffff;
  rom[28196] = 16'hffff;
  rom[28197] = 16'hffff;
  rom[28198] = 16'hffff;
  rom[28199] = 16'hffff;
  rom[28200] = 16'hffff;
  rom[28201] = 16'hffff;
  rom[28202] = 16'hffff;
  rom[28203] = 16'hffff;
  rom[28204] = 16'hffff;
  rom[28205] = 16'hffff;
  rom[28206] = 16'hffff;
  rom[28207] = 16'hffff;
  rom[28208] = 16'hffff;
  rom[28209] = 16'hffff;
  rom[28210] = 16'hff3c;
  rom[28211] = 16'hdc2f;
  rom[28212] = 16'hd269;
  rom[28213] = 16'hea07;
  rom[28214] = 16'hf227;
  rom[28215] = 16'hf206;
  rom[28216] = 16'hf227;
  rom[28217] = 16'hf227;
  rom[28218] = 16'hea27;
  rom[28219] = 16'hea26;
  rom[28220] = 16'hf226;
  rom[28221] = 16'hf207;
  rom[28222] = 16'hf228;
  rom[28223] = 16'hea06;
  rom[28224] = 16'hea26;
  rom[28225] = 16'hea06;
  rom[28226] = 16'hea27;
  rom[28227] = 16'hea06;
  rom[28228] = 16'hea26;
  rom[28229] = 16'hea06;
  rom[28230] = 16'hea27;
  rom[28231] = 16'hea26;
  rom[28232] = 16'hea46;
  rom[28233] = 16'hf206;
  rom[28234] = 16'hf227;
  rom[28235] = 16'hf1e7;
  rom[28236] = 16'hfa28;
  rom[28237] = 16'hf1e7;
  rom[28238] = 16'hfa27;
  rom[28239] = 16'hf226;
  rom[28240] = 16'hea26;
  rom[28241] = 16'hea46;
  rom[28242] = 16'hea27;
  rom[28243] = 16'hf247;
  rom[28244] = 16'hea27;
  rom[28245] = 16'hea48;
  rom[28246] = 16'hea07;
  rom[28247] = 16'hea27;
  rom[28248] = 16'hea27;
  rom[28249] = 16'hea27;
  rom[28250] = 16'hea47;
  rom[28251] = 16'he227;
  rom[28252] = 16'hea47;
  rom[28253] = 16'hea26;
  rom[28254] = 16'hf227;
  rom[28255] = 16'hf206;
  rom[28256] = 16'hfa06;
  rom[28257] = 16'hf9e6;
  rom[28258] = 16'hf227;
  rom[28259] = 16'hf206;
  rom[28260] = 16'hf226;
  rom[28261] = 16'hea26;
  rom[28262] = 16'hf246;
  rom[28263] = 16'hea07;
  rom[28264] = 16'he208;
  rom[28265] = 16'hca47;
  rom[28266] = 16'h89e3;
  rom[28267] = 16'h8304;
  rom[28268] = 16'hee90;
  rom[28269] = 16'hddcc;
  rom[28270] = 16'hd509;
  rom[28271] = 16'hb3e6;
  rom[28272] = 16'h9ae3;
  rom[28273] = 16'h8a01;
  rom[28274] = 16'h89e2;
  rom[28275] = 16'h91c2;
  rom[28276] = 16'ha1e3;
  rom[28277] = 16'hba25;
  rom[28278] = 16'hd288;
  rom[28279] = 16'hda88;
  rom[28280] = 16'hd268;
  rom[28281] = 16'hca88;
  rom[28282] = 16'hc2ca;
  rom[28283] = 16'h91a5;
  rom[28284] = 16'ha1a5;
  rom[28285] = 16'hd268;
  rom[28286] = 16'he329;
  rom[28287] = 16'hfc2b;
  rom[28288] = 16'he346;
  rom[28289] = 16'hf387;
  rom[28290] = 16'hfc2a;
  rom[28291] = 16'hfc09;
  rom[28292] = 16'hf3c9;
  rom[28293] = 16'hec28;
  rom[28294] = 16'hfe09;
  rom[28295] = 16'hff47;
  rom[28296] = 16'hffc4;
  rom[28297] = 16'hff83;
  rom[28298] = 16'hff27;
  rom[28299] = 16'hf5a7;
  rom[28300] = 16'hebe8;
  rom[28301] = 16'hf3c9;
  rom[28302] = 16'hfbc9;
  rom[28303] = 16'hfba8;
  rom[28304] = 16'hfb87;
  rom[28305] = 16'he346;
  rom[28306] = 16'hfc6c;
  rom[28307] = 16'hda87;
  rom[28308] = 16'hca49;
  rom[28309] = 16'h9925;
  rom[28310] = 16'hb146;
  rom[28311] = 16'hda48;
  rom[28312] = 16'he268;
  rom[28313] = 16'hda67;
  rom[28314] = 16'he267;
  rom[28315] = 16'he247;
  rom[28316] = 16'he247;
  rom[28317] = 16'he247;
  rom[28318] = 16'he267;
  rom[28319] = 16'hda46;
  rom[28320] = 16'hda06;
  rom[28321] = 16'hda26;
  rom[28322] = 16'he267;
  rom[28323] = 16'hda67;
  rom[28324] = 16'hd267;
  rom[28325] = 16'haa86;
  rom[28326] = 16'h7102;
  rom[28327] = 16'h9964;
  rom[28328] = 16'hda69;
  rom[28329] = 16'hea08;
  rom[28330] = 16'hf207;
  rom[28331] = 16'hea46;
  rom[28332] = 16'hea46;
  rom[28333] = 16'hf206;
  rom[28334] = 16'hf227;
  rom[28335] = 16'hea08;
  rom[28336] = 16'hf228;
  rom[28337] = 16'hf206;
  rom[28338] = 16'hf227;
  rom[28339] = 16'hf207;
  rom[28340] = 16'hf227;
  rom[28341] = 16'hea27;
  rom[28342] = 16'hda89;
  rom[28343] = 16'h8921;
  rom[28344] = 16'hab88;
  rom[28345] = 16'hf64f;
  rom[28346] = 16'hee6d;
  rom[28347] = 16'hf6cb;
  rom[28348] = 16'hff4c;
  rom[28349] = 16'hff2b;
  rom[28350] = 16'hf72a;
  rom[28351] = 16'hf729;
  rom[28352] = 16'hff49;
  rom[28353] = 16'hff48;
  rom[28354] = 16'hff28;
  rom[28355] = 16'hff28;
  rom[28356] = 16'hff29;
  rom[28357] = 16'hff29;
  rom[28358] = 16'hf72a;
  rom[28359] = 16'hf729;
  rom[28360] = 16'hf709;
  rom[28361] = 16'hff09;
  rom[28362] = 16'hff28;
  rom[28363] = 16'hf769;
  rom[28364] = 16'hf72a;
  rom[28365] = 16'hedea;
  rom[28366] = 16'h99e2;
  rom[28367] = 16'hb1e4;
  rom[28368] = 16'hd28a;
  rom[28369] = 16'hc289;
  rom[28370] = 16'hecd3;
  rom[28371] = 16'hff3c;
  rom[28372] = 16'hffbe;
  rom[28373] = 16'hfffe;
  rom[28374] = 16'hffff;
  rom[28375] = 16'hffff;
  rom[28376] = 16'hffff;
  rom[28377] = 16'hffff;
  rom[28378] = 16'hffff;
  rom[28379] = 16'hffff;
  rom[28380] = 16'hffff;
  rom[28381] = 16'hffff;
  rom[28382] = 16'hffff;
  rom[28383] = 16'hffff;
  rom[28384] = 16'hffff;
  rom[28385] = 16'hffff;
  rom[28386] = 16'hffff;
  rom[28387] = 16'hffff;
  rom[28388] = 16'hffff;
  rom[28389] = 16'hffff;
  rom[28390] = 16'hffff;
  rom[28391] = 16'hffff;
  rom[28392] = 16'hffff;
  rom[28393] = 16'hffff;
  rom[28394] = 16'hffff;
  rom[28395] = 16'hffff;
  rom[28396] = 16'hffff;
  rom[28397] = 16'hffff;
  rom[28398] = 16'hffff;
  rom[28399] = 16'hffff;
  rom[28400] = 16'hffff;
  rom[28401] = 16'hffff;
  rom[28402] = 16'hffff;
  rom[28403] = 16'hffff;
  rom[28404] = 16'hffff;
  rom[28405] = 16'hffff;
  rom[28406] = 16'hffff;
  rom[28407] = 16'hffff;
  rom[28408] = 16'hffdf;
  rom[28409] = 16'hffff;
  rom[28410] = 16'hff9d;
  rom[28411] = 16'hdcf2;
  rom[28412] = 16'hca89;
  rom[28413] = 16'hea48;
  rom[28414] = 16'hea27;
  rom[28415] = 16'hea06;
  rom[28416] = 16'he9e6;
  rom[28417] = 16'hf1e7;
  rom[28418] = 16'hea26;
  rom[28419] = 16'hf226;
  rom[28420] = 16'hf206;
  rom[28421] = 16'hf207;
  rom[28422] = 16'hea07;
  rom[28423] = 16'hea27;
  rom[28424] = 16'hea26;
  rom[28425] = 16'hea26;
  rom[28426] = 16'he206;
  rom[28427] = 16'hea06;
  rom[28428] = 16'hea06;
  rom[28429] = 16'hea06;
  rom[28430] = 16'he206;
  rom[28431] = 16'hea26;
  rom[28432] = 16'hea06;
  rom[28433] = 16'hea26;
  rom[28434] = 16'hea26;
  rom[28435] = 16'hea06;
  rom[28436] = 16'hf227;
  rom[28437] = 16'hf228;
  rom[28438] = 16'he1e6;
  rom[28439] = 16'hea27;
  rom[28440] = 16'he246;
  rom[28441] = 16'he247;
  rom[28442] = 16'hda47;
  rom[28443] = 16'he228;
  rom[28444] = 16'he208;
  rom[28445] = 16'hf229;
  rom[28446] = 16'hea07;
  rom[28447] = 16'hf228;
  rom[28448] = 16'he9e7;
  rom[28449] = 16'hf227;
  rom[28450] = 16'he1e6;
  rom[28451] = 16'hea27;
  rom[28452] = 16'hea26;
  rom[28453] = 16'hea26;
  rom[28454] = 16'hea06;
  rom[28455] = 16'hf207;
  rom[28456] = 16'hf1e6;
  rom[28457] = 16'hf206;
  rom[28458] = 16'hea06;
  rom[28459] = 16'hf226;
  rom[28460] = 16'hf206;
  rom[28461] = 16'hea26;
  rom[28462] = 16'hea26;
  rom[28463] = 16'hea07;
  rom[28464] = 16'hea07;
  rom[28465] = 16'hda89;
  rom[28466] = 16'h91e4;
  rom[28467] = 16'h6982;
  rom[28468] = 16'h9325;
  rom[28469] = 16'h8a63;
  rom[28470] = 16'h89e1;
  rom[28471] = 16'h99e2;
  rom[28472] = 16'haa04;
  rom[28473] = 16'hc246;
  rom[28474] = 16'hc266;
  rom[28475] = 16'hd287;
  rom[28476] = 16'hd246;
  rom[28477] = 16'he247;
  rom[28478] = 16'hea27;
  rom[28479] = 16'hea28;
  rom[28480] = 16'hea07;
  rom[28481] = 16'hea28;
  rom[28482] = 16'hca07;
  rom[28483] = 16'h9963;
  rom[28484] = 16'ha9a4;
  rom[28485] = 16'hda87;
  rom[28486] = 16'hfbcb;
  rom[28487] = 16'hf3ca;
  rom[28488] = 16'hca44;
  rom[28489] = 16'hf287;
  rom[28490] = 16'he245;
  rom[28491] = 16'heb07;
  rom[28492] = 16'he3a7;
  rom[28493] = 16'hfdca;
  rom[28494] = 16'hff08;
  rom[28495] = 16'hff84;
  rom[28496] = 16'hffc1;
  rom[28497] = 16'hf781;
  rom[28498] = 16'hff64;
  rom[28499] = 16'hfee9;
  rom[28500] = 16'hfd29;
  rom[28501] = 16'he3a8;
  rom[28502] = 16'he2e6;
  rom[28503] = 16'hea65;
  rom[28504] = 16'hda64;
  rom[28505] = 16'hca63;
  rom[28506] = 16'hec29;
  rom[28507] = 16'he369;
  rom[28508] = 16'hca67;
  rom[28509] = 16'ha986;
  rom[28510] = 16'hb0e4;
  rom[28511] = 16'he208;
  rom[28512] = 16'hea06;
  rom[28513] = 16'hea26;
  rom[28514] = 16'hea46;
  rom[28515] = 16'hea26;
  rom[28516] = 16'hea45;
  rom[28517] = 16'hf246;
  rom[28518] = 16'he205;
  rom[28519] = 16'hea47;
  rom[28520] = 16'he206;
  rom[28521] = 16'hea27;
  rom[28522] = 16'he206;
  rom[28523] = 16'hea47;
  rom[28524] = 16'he228;
  rom[28525] = 16'hb207;
  rom[28526] = 16'h68c0;
  rom[28527] = 16'hb1e6;
  rom[28528] = 16'hda48;
  rom[28529] = 16'he207;
  rom[28530] = 16'hf226;
  rom[28531] = 16'he205;
  rom[28532] = 16'hea25;
  rom[28533] = 16'hf206;
  rom[28534] = 16'hea06;
  rom[28535] = 16'hf208;
  rom[28536] = 16'hf208;
  rom[28537] = 16'hf207;
  rom[28538] = 16'hea06;
  rom[28539] = 16'hea07;
  rom[28540] = 16'hea07;
  rom[28541] = 16'hea07;
  rom[28542] = 16'hda68;
  rom[28543] = 16'ha984;
  rom[28544] = 16'h7962;
  rom[28545] = 16'h92e4;
  rom[28546] = 16'ha384;
  rom[28547] = 16'hb3e6;
  rom[28548] = 16'hd529;
  rom[28549] = 16'hee6c;
  rom[28550] = 16'hf70c;
  rom[28551] = 16'hff2b;
  rom[28552] = 16'hf709;
  rom[28553] = 16'hff49;
  rom[28554] = 16'hf707;
  rom[28555] = 16'hff28;
  rom[28556] = 16'hff09;
  rom[28557] = 16'hff29;
  rom[28558] = 16'hef29;
  rom[28559] = 16'hf72a;
  rom[28560] = 16'hf729;
  rom[28561] = 16'hff29;
  rom[28562] = 16'hf728;
  rom[28563] = 16'hf729;
  rom[28564] = 16'hef0b;
  rom[28565] = 16'hcce9;
  rom[28566] = 16'h8980;
  rom[28567] = 16'hc288;
  rom[28568] = 16'hc2ca;
  rom[28569] = 16'hdc91;
  rom[28570] = 16'hfeda;
  rom[28571] = 16'hffbe;
  rom[28572] = 16'hffff;
  rom[28573] = 16'hffff;
  rom[28574] = 16'hffff;
  rom[28575] = 16'hffff;
  rom[28576] = 16'hffff;
  rom[28577] = 16'hffff;
  rom[28578] = 16'hffff;
  rom[28579] = 16'hffff;
  rom[28580] = 16'hffff;
  rom[28581] = 16'hffff;
  rom[28582] = 16'hffff;
  rom[28583] = 16'hffff;
  rom[28584] = 16'hffff;
  rom[28585] = 16'hffff;
  rom[28586] = 16'hffff;
  rom[28587] = 16'hffff;
  rom[28588] = 16'hffff;
  rom[28589] = 16'hffff;
  rom[28590] = 16'hffff;
  rom[28591] = 16'hffff;
  rom[28592] = 16'hffff;
  rom[28593] = 16'hffff;
  rom[28594] = 16'hffff;
  rom[28595] = 16'hffff;
  rom[28596] = 16'hffff;
  rom[28597] = 16'hffff;
  rom[28598] = 16'hffff;
  rom[28599] = 16'hffff;
  rom[28600] = 16'hffff;
  rom[28601] = 16'hffff;
  rom[28602] = 16'hffff;
  rom[28603] = 16'hffff;
  rom[28604] = 16'hffff;
  rom[28605] = 16'hffff;
  rom[28606] = 16'hffff;
  rom[28607] = 16'hffff;
  rom[28608] = 16'hffff;
  rom[28609] = 16'hffff;
  rom[28610] = 16'hffbe;
  rom[28611] = 16'hfe99;
  rom[28612] = 16'hb289;
  rom[28613] = 16'hda07;
  rom[28614] = 16'hfa68;
  rom[28615] = 16'hf1e6;
  rom[28616] = 16'hfa89;
  rom[28617] = 16'he9e6;
  rom[28618] = 16'hf247;
  rom[28619] = 16'hea05;
  rom[28620] = 16'hf227;
  rom[28621] = 16'hf227;
  rom[28622] = 16'hea27;
  rom[28623] = 16'hea26;
  rom[28624] = 16'hea47;
  rom[28625] = 16'hea26;
  rom[28626] = 16'hea26;
  rom[28627] = 16'hea06;
  rom[28628] = 16'hea27;
  rom[28629] = 16'hea06;
  rom[28630] = 16'hea26;
  rom[28631] = 16'hea06;
  rom[28632] = 16'hea27;
  rom[28633] = 16'hea26;
  rom[28634] = 16'hea26;
  rom[28635] = 16'hea26;
  rom[28636] = 16'he1e7;
  rom[28637] = 16'he207;
  rom[28638] = 16'he249;
  rom[28639] = 16'hd227;
  rom[28640] = 16'hdaa8;
  rom[28641] = 16'hd287;
  rom[28642] = 16'hd247;
  rom[28643] = 16'hd247;
  rom[28644] = 16'he269;
  rom[28645] = 16'hd9e7;
  rom[28646] = 16'hf249;
  rom[28647] = 16'he186;
  rom[28648] = 16'hfa09;
  rom[28649] = 16'hf1e7;
  rom[28650] = 16'hfa27;
  rom[28651] = 16'hf206;
  rom[28652] = 16'hf247;
  rom[28653] = 16'hea06;
  rom[28654] = 16'hf226;
  rom[28655] = 16'hf227;
  rom[28656] = 16'hf227;
  rom[28657] = 16'hf207;
  rom[28658] = 16'hea47;
  rom[28659] = 16'hea26;
  rom[28660] = 16'hf246;
  rom[28661] = 16'hea26;
  rom[28662] = 16'hf227;
  rom[28663] = 16'hea07;
  rom[28664] = 16'hf1e7;
  rom[28665] = 16'hea89;
  rom[28666] = 16'hb246;
  rom[28667] = 16'h5080;
  rom[28668] = 16'h81a3;
  rom[28669] = 16'hb2c7;
  rom[28670] = 16'hc2a7;
  rom[28671] = 16'hdac8;
  rom[28672] = 16'he288;
  rom[28673] = 16'hda48;
  rom[28674] = 16'he247;
  rom[28675] = 16'he226;
  rom[28676] = 16'hea47;
  rom[28677] = 16'hf226;
  rom[28678] = 16'hfa26;
  rom[28679] = 16'he985;
  rom[28680] = 16'hf9c7;
  rom[28681] = 16'hfa27;
  rom[28682] = 16'he247;
  rom[28683] = 16'h9941;
  rom[28684] = 16'ha9a3;
  rom[28685] = 16'hda66;
  rom[28686] = 16'he307;
  rom[28687] = 16'hf3ea;
  rom[28688] = 16'heb08;
  rom[28689] = 16'he9e5;
  rom[28690] = 16'hea26;
  rom[28691] = 16'he2a5;
  rom[28692] = 16'he406;
  rom[28693] = 16'hfec9;
  rom[28694] = 16'hffc7;
  rom[28695] = 16'hffa2;
  rom[28696] = 16'hffc1;
  rom[28697] = 16'hffc2;
  rom[28698] = 16'hffc4;
  rom[28699] = 16'hff47;
  rom[28700] = 16'hfe2a;
  rom[28701] = 16'hd3a4;
  rom[28702] = 16'hdac6;
  rom[28703] = 16'he205;
  rom[28704] = 16'he266;
  rom[28705] = 16'he327;
  rom[28706] = 16'hfccc;
  rom[28707] = 16'hc264;
  rom[28708] = 16'hd2c8;
  rom[28709] = 16'ha185;
  rom[28710] = 16'ha8a3;
  rom[28711] = 16'hea69;
  rom[28712] = 16'he1c6;
  rom[28713] = 16'hea25;
  rom[28714] = 16'hf266;
  rom[28715] = 16'hea25;
  rom[28716] = 16'hea26;
  rom[28717] = 16'hea05;
  rom[28718] = 16'hf246;
  rom[28719] = 16'hf226;
  rom[28720] = 16'hea47;
  rom[28721] = 16'hf247;
  rom[28722] = 16'hf247;
  rom[28723] = 16'hea07;
  rom[28724] = 16'he208;
  rom[28725] = 16'hb1c6;
  rom[28726] = 16'h6041;
  rom[28727] = 16'hb1e5;
  rom[28728] = 16'hea49;
  rom[28729] = 16'hf228;
  rom[28730] = 16'hf227;
  rom[28731] = 16'hea45;
  rom[28732] = 16'hf226;
  rom[28733] = 16'hf1e6;
  rom[28734] = 16'hf227;
  rom[28735] = 16'hea07;
  rom[28736] = 16'hf227;
  rom[28737] = 16'hf206;
  rom[28738] = 16'hea46;
  rom[28739] = 16'hea26;
  rom[28740] = 16'hea28;
  rom[28741] = 16'hf227;
  rom[28742] = 16'he207;
  rom[28743] = 16'hd247;
  rom[28744] = 16'hb225;
  rom[28745] = 16'h99e2;
  rom[28746] = 16'h91c1;
  rom[28747] = 16'h8180;
  rom[28748] = 16'h7121;
  rom[28749] = 16'h9303;
  rom[28750] = 16'he60b;
  rom[28751] = 16'hff0d;
  rom[28752] = 16'hf70b;
  rom[28753] = 16'hff2a;
  rom[28754] = 16'hff0a;
  rom[28755] = 16'hff29;
  rom[28756] = 16'hff2a;
  rom[28757] = 16'hff29;
  rom[28758] = 16'hf74a;
  rom[28759] = 16'hffab;
  rom[28760] = 16'he687;
  rom[28761] = 16'hff09;
  rom[28762] = 16'hf6e8;
  rom[28763] = 16'hef2b;
  rom[28764] = 16'hf72e;
  rom[28765] = 16'h9b45;
  rom[28766] = 16'h9204;
  rom[28767] = 16'hc30a;
  rom[28768] = 16'he4d2;
  rom[28769] = 16'hfeda;
  rom[28770] = 16'hfffe;
  rom[28771] = 16'hffff;
  rom[28772] = 16'hffff;
  rom[28773] = 16'hffff;
  rom[28774] = 16'hffff;
  rom[28775] = 16'hffff;
  rom[28776] = 16'hffff;
  rom[28777] = 16'hffff;
  rom[28778] = 16'hffff;
  rom[28779] = 16'hffff;
  rom[28780] = 16'hffff;
  rom[28781] = 16'hffff;
  rom[28782] = 16'hffff;
  rom[28783] = 16'hffff;
  rom[28784] = 16'hffff;
  rom[28785] = 16'hffff;
  rom[28786] = 16'hffff;
  rom[28787] = 16'hffff;
  rom[28788] = 16'hffff;
  rom[28789] = 16'hffff;
  rom[28790] = 16'hffff;
  rom[28791] = 16'hffff;
  rom[28792] = 16'hffff;
  rom[28793] = 16'hffff;
  rom[28794] = 16'hffff;
  rom[28795] = 16'hffff;
  rom[28796] = 16'hffff;
  rom[28797] = 16'hffff;
  rom[28798] = 16'hffff;
  rom[28799] = 16'hffff;
  rom[28800] = 16'hffff;
  rom[28801] = 16'hffff;
  rom[28802] = 16'hffff;
  rom[28803] = 16'hffff;
  rom[28804] = 16'hffff;
  rom[28805] = 16'hffff;
  rom[28806] = 16'hffff;
  rom[28807] = 16'hffff;
  rom[28808] = 16'hffff;
  rom[28809] = 16'hffff;
  rom[28810] = 16'hffde;
  rom[28811] = 16'hfefb;
  rom[28812] = 16'hc36c;
  rom[28813] = 16'hda68;
  rom[28814] = 16'hea27;
  rom[28815] = 16'hf227;
  rom[28816] = 16'hf227;
  rom[28817] = 16'he9e6;
  rom[28818] = 16'hf226;
  rom[28819] = 16'hf205;
  rom[28820] = 16'hea06;
  rom[28821] = 16'hf227;
  rom[28822] = 16'hea07;
  rom[28823] = 16'hea27;
  rom[28824] = 16'he226;
  rom[28825] = 16'hea26;
  rom[28826] = 16'hea26;
  rom[28827] = 16'hea26;
  rom[28828] = 16'he206;
  rom[28829] = 16'hea06;
  rom[28830] = 16'hea06;
  rom[28831] = 16'hea06;
  rom[28832] = 16'he206;
  rom[28833] = 16'hea26;
  rom[28834] = 16'hea26;
  rom[28835] = 16'he205;
  rom[28836] = 16'hf288;
  rom[28837] = 16'he227;
  rom[28838] = 16'hca47;
  rom[28839] = 16'hca66;
  rom[28840] = 16'h99c2;
  rom[28841] = 16'h91c2;
  rom[28842] = 16'h9a23;
  rom[28843] = 16'h9180;
  rom[28844] = 16'ha1c3;
  rom[28845] = 16'hca87;
  rom[28846] = 16'hd247;
  rom[28847] = 16'he248;
  rom[28848] = 16'hea07;
  rom[28849] = 16'hfa07;
  rom[28850] = 16'hf1c6;
  rom[28851] = 16'hfa07;
  rom[28852] = 16'hf206;
  rom[28853] = 16'hea26;
  rom[28854] = 16'hea06;
  rom[28855] = 16'hea27;
  rom[28856] = 16'hea07;
  rom[28857] = 16'hea07;
  rom[28858] = 16'hea27;
  rom[28859] = 16'hea27;
  rom[28860] = 16'hea25;
  rom[28861] = 16'hf226;
  rom[28862] = 16'hea06;
  rom[28863] = 16'hfa28;
  rom[28864] = 16'he985;
  rom[28865] = 16'hea07;
  rom[28866] = 16'hba67;
  rom[28867] = 16'h68a0;
  rom[28868] = 16'h91c5;
  rom[28869] = 16'hc268;
  rom[28870] = 16'hd247;
  rom[28871] = 16'he227;
  rom[28872] = 16'hea07;
  rom[28873] = 16'hf207;
  rom[28874] = 16'he9e6;
  rom[28875] = 16'hf227;
  rom[28876] = 16'he9e5;
  rom[28877] = 16'hf206;
  rom[28878] = 16'hf1e6;
  rom[28879] = 16'hfa07;
  rom[28880] = 16'hf1e6;
  rom[28881] = 16'hf226;
  rom[28882] = 16'hd225;
  rom[28883] = 16'ha1a3;
  rom[28884] = 16'ha162;
  rom[28885] = 16'hda46;
  rom[28886] = 16'hda86;
  rom[28887] = 16'hfbaa;
  rom[28888] = 16'heb08;
  rom[28889] = 16'hea26;
  rom[28890] = 16'he245;
  rom[28891] = 16'hdae4;
  rom[28892] = 16'hf547;
  rom[28893] = 16'hff88;
  rom[28894] = 16'hff83;
  rom[28895] = 16'hffc2;
  rom[28896] = 16'hff61;
  rom[28897] = 16'hff82;
  rom[28898] = 16'hff62;
  rom[28899] = 16'hff85;
  rom[28900] = 16'hfee7;
  rom[28901] = 16'hf527;
  rom[28902] = 16'hcae3;
  rom[28903] = 16'he265;
  rom[28904] = 16'hda24;
  rom[28905] = 16'hfc2c;
  rom[28906] = 16'he368;
  rom[28907] = 16'heb08;
  rom[28908] = 16'hba05;
  rom[28909] = 16'h9984;
  rom[28910] = 16'ha144;
  rom[28911] = 16'hda68;
  rom[28912] = 16'hda26;
  rom[28913] = 16'he267;
  rom[28914] = 16'hda25;
  rom[28915] = 16'he246;
  rom[28916] = 16'he246;
  rom[28917] = 16'he246;
  rom[28918] = 16'he226;
  rom[28919] = 16'hea27;
  rom[28920] = 16'he247;
  rom[28921] = 16'he227;
  rom[28922] = 16'hda07;
  rom[28923] = 16'hea69;
  rom[28924] = 16'hda28;
  rom[28925] = 16'ha1c6;
  rom[28926] = 16'h68a0;
  rom[28927] = 16'hc227;
  rom[28928] = 16'he1e7;
  rom[28929] = 16'hfa29;
  rom[28930] = 16'hea06;
  rom[28931] = 16'hea26;
  rom[28932] = 16'hea26;
  rom[28933] = 16'hf1e7;
  rom[28934] = 16'hf207;
  rom[28935] = 16'hf207;
  rom[28936] = 16'hea07;
  rom[28937] = 16'hf226;
  rom[28938] = 16'hea26;
  rom[28939] = 16'hea27;
  rom[28940] = 16'he207;
  rom[28941] = 16'hf207;
  rom[28942] = 16'hea07;
  rom[28943] = 16'hea48;
  rom[28944] = 16'hd247;
  rom[28945] = 16'hca66;
  rom[28946] = 16'hca86;
  rom[28947] = 16'hca87;
  rom[28948] = 16'hb245;
  rom[28949] = 16'h81e1;
  rom[28950] = 16'h7a61;
  rom[28951] = 16'he5ec;
  rom[28952] = 16'heecc;
  rom[28953] = 16'hff4c;
  rom[28954] = 16'hff0a;
  rom[28955] = 16'hff29;
  rom[28956] = 16'hf708;
  rom[28957] = 16'hff29;
  rom[28958] = 16'hf728;
  rom[28959] = 16'hf729;
  rom[28960] = 16'hff4a;
  rom[28961] = 16'hfee8;
  rom[28962] = 16'hf6e9;
  rom[28963] = 16'hf72d;
  rom[28964] = 16'hbdcc;
  rom[28965] = 16'h6223;
  rom[28966] = 16'h9b4a;
  rom[28967] = 16'hed55;
  rom[28968] = 16'hfeda;
  rom[28969] = 16'hffde;
  rom[28970] = 16'hfffe;
  rom[28971] = 16'hffff;
  rom[28972] = 16'hffff;
  rom[28973] = 16'hffff;
  rom[28974] = 16'hffff;
  rom[28975] = 16'hffff;
  rom[28976] = 16'hffff;
  rom[28977] = 16'hffff;
  rom[28978] = 16'hffff;
  rom[28979] = 16'hffff;
  rom[28980] = 16'hffff;
  rom[28981] = 16'hffff;
  rom[28982] = 16'hffff;
  rom[28983] = 16'hffff;
  rom[28984] = 16'hffff;
  rom[28985] = 16'hffff;
  rom[28986] = 16'hffff;
  rom[28987] = 16'hffff;
  rom[28988] = 16'hffff;
  rom[28989] = 16'hffff;
  rom[28990] = 16'hffff;
  rom[28991] = 16'hffff;
  rom[28992] = 16'hffff;
  rom[28993] = 16'hffff;
  rom[28994] = 16'hffff;
  rom[28995] = 16'hffff;
  rom[28996] = 16'hffff;
  rom[28997] = 16'hffff;
  rom[28998] = 16'hffff;
  rom[28999] = 16'hffff;
  rom[29000] = 16'hffff;
  rom[29001] = 16'hffff;
  rom[29002] = 16'hffff;
  rom[29003] = 16'hffff;
  rom[29004] = 16'hffff;
  rom[29005] = 16'hffff;
  rom[29006] = 16'hffff;
  rom[29007] = 16'hffff;
  rom[29008] = 16'hffff;
  rom[29009] = 16'hffff;
  rom[29010] = 16'hffff;
  rom[29011] = 16'hff9d;
  rom[29012] = 16'hf533;
  rom[29013] = 16'hca68;
  rom[29014] = 16'hf269;
  rom[29015] = 16'he1c6;
  rom[29016] = 16'hf227;
  rom[29017] = 16'hf207;
  rom[29018] = 16'hf227;
  rom[29019] = 16'hf226;
  rom[29020] = 16'hf226;
  rom[29021] = 16'hea27;
  rom[29022] = 16'hea48;
  rom[29023] = 16'hea26;
  rom[29024] = 16'hea46;
  rom[29025] = 16'hea26;
  rom[29026] = 16'hea47;
  rom[29027] = 16'hea26;
  rom[29028] = 16'hea26;
  rom[29029] = 16'hea06;
  rom[29030] = 16'hea27;
  rom[29031] = 16'hea06;
  rom[29032] = 16'hf226;
  rom[29033] = 16'hf206;
  rom[29034] = 16'hfa26;
  rom[29035] = 16'hf227;
  rom[29036] = 16'hea27;
  rom[29037] = 16'hda47;
  rom[29038] = 16'hd2a7;
  rom[29039] = 16'h99e3;
  rom[29040] = 16'ha2c3;
  rom[29041] = 16'hdd2b;
  rom[29042] = 16'hf5cd;
  rom[29043] = 16'he58c;
  rom[29044] = 16'h92c2;
  rom[29045] = 16'h7980;
  rom[29046] = 16'haa24;
  rom[29047] = 16'hca86;
  rom[29048] = 16'he247;
  rom[29049] = 16'he9e5;
  rom[29050] = 16'hf9e7;
  rom[29051] = 16'hf1e6;
  rom[29052] = 16'hf206;
  rom[29053] = 16'hea27;
  rom[29054] = 16'hea47;
  rom[29055] = 16'hea27;
  rom[29056] = 16'hf227;
  rom[29057] = 16'hf207;
  rom[29058] = 16'hea48;
  rom[29059] = 16'hea26;
  rom[29060] = 16'hf245;
  rom[29061] = 16'hf225;
  rom[29062] = 16'hf248;
  rom[29063] = 16'he9c6;
  rom[29064] = 16'hfa07;
  rom[29065] = 16'hea48;
  rom[29066] = 16'hc288;
  rom[29067] = 16'h7902;
  rom[29068] = 16'h9985;
  rom[29069] = 16'hca68;
  rom[29070] = 16'he268;
  rom[29071] = 16'hea07;
  rom[29072] = 16'hfa07;
  rom[29073] = 16'hf1e7;
  rom[29074] = 16'hf1e7;
  rom[29075] = 16'hea06;
  rom[29076] = 16'hea27;
  rom[29077] = 16'hea47;
  rom[29078] = 16'hf228;
  rom[29079] = 16'he228;
  rom[29080] = 16'he207;
  rom[29081] = 16'hea47;
  rom[29082] = 16'hdaa8;
  rom[29083] = 16'haa25;
  rom[29084] = 16'h9943;
  rom[29085] = 16'hd206;
  rom[29086] = 16'hda46;
  rom[29087] = 16'hf368;
  rom[29088] = 16'hfc2b;
  rom[29089] = 16'heae8;
  rom[29090] = 16'hd265;
  rom[29091] = 16'he407;
  rom[29092] = 16'hfe8a;
  rom[29093] = 16'hff86;
  rom[29094] = 16'hff82;
  rom[29095] = 16'hffa3;
  rom[29096] = 16'hff23;
  rom[29097] = 16'hff23;
  rom[29098] = 16'hff22;
  rom[29099] = 16'hff84;
  rom[29100] = 16'hff26;
  rom[29101] = 16'hfe28;
  rom[29102] = 16'hdba4;
  rom[29103] = 16'he2a4;
  rom[29104] = 16'hf348;
  rom[29105] = 16'hfcae;
  rom[29106] = 16'hdae8;
  rom[29107] = 16'hda47;
  rom[29108] = 16'hd2c9;
  rom[29109] = 16'h8122;
  rom[29110] = 16'haa26;
  rom[29111] = 16'hc267;
  rom[29112] = 16'hcaa8;
  rom[29113] = 16'hcaa7;
  rom[29114] = 16'hcac7;
  rom[29115] = 16'hcac7;
  rom[29116] = 16'hcaa7;
  rom[29117] = 16'hca87;
  rom[29118] = 16'hd2c8;
  rom[29119] = 16'hca87;
  rom[29120] = 16'hd2a8;
  rom[29121] = 16'hca88;
  rom[29122] = 16'hd2a9;
  rom[29123] = 16'hca68;
  rom[29124] = 16'hc248;
  rom[29125] = 16'h8944;
  rom[29126] = 16'h7943;
  rom[29127] = 16'hd269;
  rom[29128] = 16'hf1e8;
  rom[29129] = 16'hfa09;
  rom[29130] = 16'hea07;
  rom[29131] = 16'he226;
  rom[29132] = 16'hea47;
  rom[29133] = 16'hf208;
  rom[29134] = 16'hf228;
  rom[29135] = 16'hf207;
  rom[29136] = 16'hf226;
  rom[29137] = 16'hf225;
  rom[29138] = 16'hea66;
  rom[29139] = 16'hea46;
  rom[29140] = 16'hea47;
  rom[29141] = 16'hf207;
  rom[29142] = 16'hf1a7;
  rom[29143] = 16'hf1e7;
  rom[29144] = 16'hea28;
  rom[29145] = 16'hda26;
  rom[29146] = 16'he247;
  rom[29147] = 16'hda28;
  rom[29148] = 16'hca47;
  rom[29149] = 16'hb2c6;
  rom[29150] = 16'h7160;
  rom[29151] = 16'ha3c5;
  rom[29152] = 16'hf6ad;
  rom[29153] = 16'hff2d;
  rom[29154] = 16'hff2a;
  rom[29155] = 16'hff28;
  rom[29156] = 16'hff49;
  rom[29157] = 16'hff27;
  rom[29158] = 16'hff49;
  rom[29159] = 16'hff6a;
  rom[29160] = 16'heee8;
  rom[29161] = 16'hff29;
  rom[29162] = 16'hf688;
  rom[29163] = 16'he6cd;
  rom[29164] = 16'h73a5;
  rom[29165] = 16'h7b6a;
  rom[29166] = 16'hf699;
  rom[29167] = 16'hff5d;
  rom[29168] = 16'hff9e;
  rom[29169] = 16'hffff;
  rom[29170] = 16'hffff;
  rom[29171] = 16'hffff;
  rom[29172] = 16'hffff;
  rom[29173] = 16'hffff;
  rom[29174] = 16'hffff;
  rom[29175] = 16'hffff;
  rom[29176] = 16'hffff;
  rom[29177] = 16'hffff;
  rom[29178] = 16'hffff;
  rom[29179] = 16'hffff;
  rom[29180] = 16'hffff;
  rom[29181] = 16'hffff;
  rom[29182] = 16'hffff;
  rom[29183] = 16'hffff;
  rom[29184] = 16'hffff;
  rom[29185] = 16'hffff;
  rom[29186] = 16'hffff;
  rom[29187] = 16'hffff;
  rom[29188] = 16'hffff;
  rom[29189] = 16'hffff;
  rom[29190] = 16'hffff;
  rom[29191] = 16'hffff;
  rom[29192] = 16'hffff;
  rom[29193] = 16'hffff;
  rom[29194] = 16'hffff;
  rom[29195] = 16'hffff;
  rom[29196] = 16'hffff;
  rom[29197] = 16'hffff;
  rom[29198] = 16'hffff;
  rom[29199] = 16'hffff;
  rom[29200] = 16'hffff;
  rom[29201] = 16'hffff;
  rom[29202] = 16'hffff;
  rom[29203] = 16'hffff;
  rom[29204] = 16'hffff;
  rom[29205] = 16'hffff;
  rom[29206] = 16'hffff;
  rom[29207] = 16'hffff;
  rom[29208] = 16'hffff;
  rom[29209] = 16'hffff;
  rom[29210] = 16'hffff;
  rom[29211] = 16'hffde;
  rom[29212] = 16'hfeb9;
  rom[29213] = 16'hd30c;
  rom[29214] = 16'hda27;
  rom[29215] = 16'hf247;
  rom[29216] = 16'hea07;
  rom[29217] = 16'hf227;
  rom[29218] = 16'hea06;
  rom[29219] = 16'hf207;
  rom[29220] = 16'hf206;
  rom[29221] = 16'hea26;
  rom[29222] = 16'he226;
  rom[29223] = 16'hea26;
  rom[29224] = 16'hea26;
  rom[29225] = 16'hea27;
  rom[29226] = 16'he226;
  rom[29227] = 16'hea26;
  rom[29228] = 16'hea06;
  rom[29229] = 16'hea06;
  rom[29230] = 16'hea06;
  rom[29231] = 16'hea06;
  rom[29232] = 16'hea06;
  rom[29233] = 16'hf206;
  rom[29234] = 16'hea06;
  rom[29235] = 16'hf227;
  rom[29236] = 16'hea06;
  rom[29237] = 16'he268;
  rom[29238] = 16'hba46;
  rom[29239] = 16'h9201;
  rom[29240] = 16'hdd6c;
  rom[29241] = 16'hfeee;
  rom[29242] = 16'hf6ec;
  rom[29243] = 16'hf6cc;
  rom[29244] = 16'hf68c;
  rom[29245] = 16'hb426;
  rom[29246] = 16'h8222;
  rom[29247] = 16'ha223;
  rom[29248] = 16'hca86;
  rom[29249] = 16'he226;
  rom[29250] = 16'hea06;
  rom[29251] = 16'hf206;
  rom[29252] = 16'hf1e6;
  rom[29253] = 16'hf207;
  rom[29254] = 16'hea06;
  rom[29255] = 16'hea27;
  rom[29256] = 16'hea07;
  rom[29257] = 16'hf207;
  rom[29258] = 16'hea07;
  rom[29259] = 16'hea26;
  rom[29260] = 16'hf225;
  rom[29261] = 16'hf245;
  rom[29262] = 16'hea06;
  rom[29263] = 16'hf228;
  rom[29264] = 16'hea07;
  rom[29265] = 16'he246;
  rom[29266] = 16'hba87;
  rom[29267] = 16'h8163;
  rom[29268] = 16'h80e3;
  rom[29269] = 16'hd269;
  rom[29270] = 16'he207;
  rom[29271] = 16'hea07;
  rom[29272] = 16'hf206;
  rom[29273] = 16'hf206;
  rom[29274] = 16'he226;
  rom[29275] = 16'hea47;
  rom[29276] = 16'he227;
  rom[29277] = 16'he208;
  rom[29278] = 16'hda08;
  rom[29279] = 16'hda48;
  rom[29280] = 16'hd247;
  rom[29281] = 16'hda88;
  rom[29282] = 16'hba87;
  rom[29283] = 16'h9a25;
  rom[29284] = 16'h8102;
  rom[29285] = 16'hd247;
  rom[29286] = 16'he266;
  rom[29287] = 16'hda44;
  rom[29288] = 16'hfc2a;
  rom[29289] = 16'hf3c9;
  rom[29290] = 16'hcb46;
  rom[29291] = 16'hfded;
  rom[29292] = 16'hfeea;
  rom[29293] = 16'hff46;
  rom[29294] = 16'hff64;
  rom[29295] = 16'hff45;
  rom[29296] = 16'hfee5;
  rom[29297] = 16'hff27;
  rom[29298] = 16'hff25;
  rom[29299] = 16'hff87;
  rom[29300] = 16'hff26;
  rom[29301] = 16'hfeea;
  rom[29302] = 16'hfd49;
  rom[29303] = 16'hd324;
  rom[29304] = 16'hf42b;
  rom[29305] = 16'he2e8;
  rom[29306] = 16'hda88;
  rom[29307] = 16'hd228;
  rom[29308] = 16'hb226;
  rom[29309] = 16'h7121;
  rom[29310] = 16'h89e2;
  rom[29311] = 16'h9223;
  rom[29312] = 16'h9243;
  rom[29313] = 16'h9244;
  rom[29314] = 16'h9264;
  rom[29315] = 16'h9a64;
  rom[29316] = 16'h9263;
  rom[29317] = 16'h9263;
  rom[29318] = 16'h8a21;
  rom[29319] = 16'h8a02;
  rom[29320] = 16'h81e1;
  rom[29321] = 16'h81a1;
  rom[29322] = 16'h8a22;
  rom[29323] = 16'h89c3;
  rom[29324] = 16'h91e3;
  rom[29325] = 16'h6902;
  rom[29326] = 16'h8164;
  rom[29327] = 16'hd268;
  rom[29328] = 16'hf1e7;
  rom[29329] = 16'hf9c7;
  rom[29330] = 16'he9e7;
  rom[29331] = 16'hea48;
  rom[29332] = 16'hea27;
  rom[29333] = 16'hf228;
  rom[29334] = 16'hea06;
  rom[29335] = 16'hf226;
  rom[29336] = 16'hf206;
  rom[29337] = 16'hf225;
  rom[29338] = 16'he245;
  rom[29339] = 16'he246;
  rom[29340] = 16'he226;
  rom[29341] = 16'hfa07;
  rom[29342] = 16'hf9e6;
  rom[29343] = 16'hf9c7;
  rom[29344] = 16'he9e7;
  rom[29345] = 16'hea47;
  rom[29346] = 16'he226;
  rom[29347] = 16'hea28;
  rom[29348] = 16'hda88;
  rom[29349] = 16'hcac8;
  rom[29350] = 16'h8a43;
  rom[29351] = 16'h82c2;
  rom[29352] = 16'he66c;
  rom[29353] = 16'hf72d;
  rom[29354] = 16'hef2a;
  rom[29355] = 16'hf728;
  rom[29356] = 16'hff27;
  rom[29357] = 16'hff07;
  rom[29358] = 16'hf709;
  rom[29359] = 16'he6e8;
  rom[29360] = 16'hff6a;
  rom[29361] = 16'hf72a;
  rom[29362] = 16'hf72c;
  rom[29363] = 16'hb549;
  rom[29364] = 16'h5ae5;
  rom[29365] = 16'hd677;
  rom[29366] = 16'hffbe;
  rom[29367] = 16'hffbf;
  rom[29368] = 16'hffff;
  rom[29369] = 16'hffff;
  rom[29370] = 16'hffff;
  rom[29371] = 16'hffff;
  rom[29372] = 16'hffff;
  rom[29373] = 16'hffff;
  rom[29374] = 16'hffff;
  rom[29375] = 16'hffff;
  rom[29376] = 16'hffff;
  rom[29377] = 16'hffff;
  rom[29378] = 16'hffff;
  rom[29379] = 16'hffff;
  rom[29380] = 16'hffff;
  rom[29381] = 16'hffff;
  rom[29382] = 16'hffff;
  rom[29383] = 16'hffff;
  rom[29384] = 16'hffff;
  rom[29385] = 16'hffff;
  rom[29386] = 16'hffff;
  rom[29387] = 16'hffff;
  rom[29388] = 16'hffff;
  rom[29389] = 16'hffff;
  rom[29390] = 16'hffff;
  rom[29391] = 16'hffff;
  rom[29392] = 16'hffff;
  rom[29393] = 16'hffff;
  rom[29394] = 16'hffff;
  rom[29395] = 16'hffff;
  rom[29396] = 16'hffff;
  rom[29397] = 16'hffff;
  rom[29398] = 16'hffff;
  rom[29399] = 16'hffff;
  rom[29400] = 16'hffff;
  rom[29401] = 16'hffff;
  rom[29402] = 16'hffff;
  rom[29403] = 16'hffff;
  rom[29404] = 16'hffff;
  rom[29405] = 16'hffff;
  rom[29406] = 16'hffff;
  rom[29407] = 16'hffff;
  rom[29408] = 16'hffff;
  rom[29409] = 16'hffff;
  rom[29410] = 16'hffff;
  rom[29411] = 16'hffdf;
  rom[29412] = 16'hff7d;
  rom[29413] = 16'he450;
  rom[29414] = 16'hd267;
  rom[29415] = 16'hea47;
  rom[29416] = 16'hf247;
  rom[29417] = 16'hf227;
  rom[29418] = 16'hf207;
  rom[29419] = 16'hf207;
  rom[29420] = 16'hf227;
  rom[29421] = 16'hea26;
  rom[29422] = 16'hea46;
  rom[29423] = 16'hea27;
  rom[29424] = 16'hea48;
  rom[29425] = 16'hea27;
  rom[29426] = 16'hea27;
  rom[29427] = 16'hf206;
  rom[29428] = 16'hf227;
  rom[29429] = 16'hf206;
  rom[29430] = 16'hf226;
  rom[29431] = 16'hf206;
  rom[29432] = 16'hf227;
  rom[29433] = 16'hea07;
  rom[29434] = 16'hf227;
  rom[29435] = 16'he9e6;
  rom[29436] = 16'hf206;
  rom[29437] = 16'hda26;
  rom[29438] = 16'hc246;
  rom[29439] = 16'h9223;
  rom[29440] = 16'hee2e;
  rom[29441] = 16'heeea;
  rom[29442] = 16'hff8c;
  rom[29443] = 16'hf72a;
  rom[29444] = 16'hfeec;
  rom[29445] = 16'hf6ac;
  rom[29446] = 16'hcd09;
  rom[29447] = 16'h9261;
  rom[29448] = 16'h99e2;
  rom[29449] = 16'hca46;
  rom[29450] = 16'he247;
  rom[29451] = 16'hea46;
  rom[29452] = 16'hf247;
  rom[29453] = 16'hf227;
  rom[29454] = 16'hf207;
  rom[29455] = 16'hea47;
  rom[29456] = 16'hea27;
  rom[29457] = 16'hf207;
  rom[29458] = 16'hf227;
  rom[29459] = 16'hf225;
  rom[29460] = 16'hf245;
  rom[29461] = 16'hea46;
  rom[29462] = 16'hf227;
  rom[29463] = 16'hea07;
  rom[29464] = 16'hea88;
  rom[29465] = 16'hd2c7;
  rom[29466] = 16'h91c3;
  rom[29467] = 16'h6901;
  rom[29468] = 16'h70e3;
  rom[29469] = 16'hc228;
  rom[29470] = 16'he249;
  rom[29471] = 16'he1e7;
  rom[29472] = 16'hea47;
  rom[29473] = 16'he226;
  rom[29474] = 16'he267;
  rom[29475] = 16'he268;
  rom[29476] = 16'he2a9;
  rom[29477] = 16'hda68;
  rom[29478] = 16'hda47;
  rom[29479] = 16'hca87;
  rom[29480] = 16'hc267;
  rom[29481] = 16'ha1a4;
  rom[29482] = 16'h8183;
  rom[29483] = 16'h6141;
  rom[29484] = 16'h7121;
  rom[29485] = 16'ha9c3;
  rom[29486] = 16'he267;
  rom[29487] = 16'hda04;
  rom[29488] = 16'he2a5;
  rom[29489] = 16'hfccc;
  rom[29490] = 16'hfd2c;
  rom[29491] = 16'hfe4e;
  rom[29492] = 16'hff0c;
  rom[29493] = 16'hff29;
  rom[29494] = 16'hff08;
  rom[29495] = 16'hfec9;
  rom[29496] = 16'hfeaa;
  rom[29497] = 16'hfecb;
  rom[29498] = 16'hfeeb;
  rom[29499] = 16'hfeea;
  rom[29500] = 16'hff0b;
  rom[29501] = 16'hfecb;
  rom[29502] = 16'hfe6d;
  rom[29503] = 16'hec89;
  rom[29504] = 16'hfc2c;
  rom[29505] = 16'he289;
  rom[29506] = 16'he249;
  rom[29507] = 16'hca67;
  rom[29508] = 16'ha204;
  rom[29509] = 16'ha325;
  rom[29510] = 16'hdd6b;
  rom[29511] = 16'hee6c;
  rom[29512] = 16'hf6ac;
  rom[29513] = 16'hf64c;
  rom[29514] = 16'hf66d;
  rom[29515] = 16'hf66c;
  rom[29516] = 16'hfeee;
  rom[29517] = 16'hf68d;
  rom[29518] = 16'hee0c;
  rom[29519] = 16'hddcb;
  rom[29520] = 16'he5cc;
  rom[29521] = 16'hcd0a;
  rom[29522] = 16'hcd0b;
  rom[29523] = 16'hc4aa;
  rom[29524] = 16'hccab;
  rom[29525] = 16'h79e3;
  rom[29526] = 16'h91e5;
  rom[29527] = 16'hda69;
  rom[29528] = 16'hfa08;
  rom[29529] = 16'hf9e6;
  rom[29530] = 16'hfa08;
  rom[29531] = 16'he9e8;
  rom[29532] = 16'hea28;
  rom[29533] = 16'hea27;
  rom[29534] = 16'hea25;
  rom[29535] = 16'hf205;
  rom[29536] = 16'hfa06;
  rom[29537] = 16'hea26;
  rom[29538] = 16'hea66;
  rom[29539] = 16'he246;
  rom[29540] = 16'hea27;
  rom[29541] = 16'hf206;
  rom[29542] = 16'hfa07;
  rom[29543] = 16'hf207;
  rom[29544] = 16'hea47;
  rom[29545] = 16'hda67;
  rom[29546] = 16'hda47;
  rom[29547] = 16'hda69;
  rom[29548] = 16'hca29;
  rom[29549] = 16'hc2c9;
  rom[29550] = 16'ha2a6;
  rom[29551] = 16'h8282;
  rom[29552] = 16'hf6d0;
  rom[29553] = 16'hef0c;
  rom[29554] = 16'hf72a;
  rom[29555] = 16'hf729;
  rom[29556] = 16'hff29;
  rom[29557] = 16'hff29;
  rom[29558] = 16'hff2a;
  rom[29559] = 16'hf72b;
  rom[29560] = 16'hf72b;
  rom[29561] = 16'he6eb;
  rom[29562] = 16'hd64c;
  rom[29563] = 16'h6322;
  rom[29564] = 16'hb592;
  rom[29565] = 16'hffde;
  rom[29566] = 16'hffff;
  rom[29567] = 16'hffff;
  rom[29568] = 16'hffff;
  rom[29569] = 16'hffff;
  rom[29570] = 16'hffff;
  rom[29571] = 16'hffff;
  rom[29572] = 16'hffff;
  rom[29573] = 16'hffff;
  rom[29574] = 16'hffff;
  rom[29575] = 16'hffff;
  rom[29576] = 16'hffff;
  rom[29577] = 16'hffff;
  rom[29578] = 16'hffff;
  rom[29579] = 16'hffff;
  rom[29580] = 16'hffff;
  rom[29581] = 16'hffff;
  rom[29582] = 16'hffff;
  rom[29583] = 16'hffff;
  rom[29584] = 16'hffff;
  rom[29585] = 16'hffff;
  rom[29586] = 16'hffff;
  rom[29587] = 16'hffff;
  rom[29588] = 16'hffff;
  rom[29589] = 16'hffff;
  rom[29590] = 16'hffff;
  rom[29591] = 16'hffff;
  rom[29592] = 16'hffff;
  rom[29593] = 16'hffff;
  rom[29594] = 16'hffff;
  rom[29595] = 16'hffff;
  rom[29596] = 16'hffff;
  rom[29597] = 16'hffff;
  rom[29598] = 16'hffff;
  rom[29599] = 16'hffff;
  rom[29600] = 16'hffff;
  rom[29601] = 16'hffff;
  rom[29602] = 16'hffff;
  rom[29603] = 16'hffff;
  rom[29604] = 16'hffff;
  rom[29605] = 16'hffff;
  rom[29606] = 16'hffff;
  rom[29607] = 16'hffff;
  rom[29608] = 16'hffff;
  rom[29609] = 16'hffff;
  rom[29610] = 16'hffff;
  rom[29611] = 16'hffff;
  rom[29612] = 16'hffbc;
  rom[29613] = 16'hed53;
  rom[29614] = 16'hcac9;
  rom[29615] = 16'he268;
  rom[29616] = 16'hea06;
  rom[29617] = 16'hf206;
  rom[29618] = 16'hf207;
  rom[29619] = 16'hf227;
  rom[29620] = 16'hea06;
  rom[29621] = 16'hf247;
  rom[29622] = 16'hea06;
  rom[29623] = 16'hea07;
  rom[29624] = 16'hea07;
  rom[29625] = 16'hea07;
  rom[29626] = 16'hea07;
  rom[29627] = 16'hea06;
  rom[29628] = 16'hea06;
  rom[29629] = 16'hf206;
  rom[29630] = 16'hf206;
  rom[29631] = 16'hf206;
  rom[29632] = 16'hea06;
  rom[29633] = 16'hf206;
  rom[29634] = 16'hea27;
  rom[29635] = 16'hfa27;
  rom[29636] = 16'hea06;
  rom[29637] = 16'hea48;
  rom[29638] = 16'hcaa8;
  rom[29639] = 16'h9263;
  rom[29640] = 16'hf64d;
  rom[29641] = 16'hff4c;
  rom[29642] = 16'heec7;
  rom[29643] = 16'hff29;
  rom[29644] = 16'hff2b;
  rom[29645] = 16'hf70c;
  rom[29646] = 16'hf6ed;
  rom[29647] = 16'hc4c7;
  rom[29648] = 16'h81e0;
  rom[29649] = 16'hb265;
  rom[29650] = 16'hca67;
  rom[29651] = 16'he227;
  rom[29652] = 16'he9e6;
  rom[29653] = 16'hea06;
  rom[29654] = 16'hea05;
  rom[29655] = 16'hf246;
  rom[29656] = 16'hea26;
  rom[29657] = 16'he9e6;
  rom[29658] = 16'hf1e6;
  rom[29659] = 16'hf206;
  rom[29660] = 16'hea25;
  rom[29661] = 16'hea27;
  rom[29662] = 16'hda07;
  rom[29663] = 16'he269;
  rom[29664] = 16'hca87;
  rom[29665] = 16'h9a02;
  rom[29666] = 16'h69c1;
  rom[29667] = 16'h9b69;
  rom[29668] = 16'h6123;
  rom[29669] = 16'hba69;
  rom[29670] = 16'hd249;
  rom[29671] = 16'he229;
  rom[29672] = 16'hda67;
  rom[29673] = 16'hda87;
  rom[29674] = 16'hca66;
  rom[29675] = 16'hba47;
  rom[29676] = 16'haa46;
  rom[29677] = 16'ha245;
  rom[29678] = 16'h89a1;
  rom[29679] = 16'h8161;
  rom[29680] = 16'h7962;
  rom[29681] = 16'h81e2;
  rom[29682] = 16'hbc27;
  rom[29683] = 16'hd54c;
  rom[29684] = 16'hb427;
  rom[29685] = 16'h9202;
  rom[29686] = 16'hca25;
  rom[29687] = 16'hea87;
  rom[29688] = 16'hda25;
  rom[29689] = 16'he348;
  rom[29690] = 16'hf4ab;
  rom[29691] = 16'hc343;
  rom[29692] = 16'he4c6;
  rom[29693] = 16'hed06;
  rom[29694] = 16'hc381;
  rom[29695] = 16'hd362;
  rom[29696] = 16'hcb23;
  rom[29697] = 16'hcb24;
  rom[29698] = 16'hc322;
  rom[29699] = 16'hcbe3;
  rom[29700] = 16'hf548;
  rom[29701] = 16'hcc24;
  rom[29702] = 16'hc363;
  rom[29703] = 16'hfccb;
  rom[29704] = 16'he307;
  rom[29705] = 16'hda46;
  rom[29706] = 16'hd267;
  rom[29707] = 16'hc286;
  rom[29708] = 16'h9201;
  rom[29709] = 16'he56a;
  rom[29710] = 16'hfecc;
  rom[29711] = 16'hff0a;
  rom[29712] = 16'hf72a;
  rom[29713] = 16'hff2b;
  rom[29714] = 16'hfeeb;
  rom[29715] = 16'hff2d;
  rom[29716] = 16'heecb;
  rom[29717] = 16'hf6ed;
  rom[29718] = 16'hff0d;
  rom[29719] = 16'hf6ed;
  rom[29720] = 16'heecd;
  rom[29721] = 16'hf6ce;
  rom[29722] = 16'hff0e;
  rom[29723] = 16'hff0f;
  rom[29724] = 16'hee4e;
  rom[29725] = 16'h8a62;
  rom[29726] = 16'ha225;
  rom[29727] = 16'he268;
  rom[29728] = 16'hf1e5;
  rom[29729] = 16'hf1c6;
  rom[29730] = 16'hf207;
  rom[29731] = 16'hf228;
  rom[29732] = 16'he9e7;
  rom[29733] = 16'hea06;
  rom[29734] = 16'hf206;
  rom[29735] = 16'hf206;
  rom[29736] = 16'hf226;
  rom[29737] = 16'hf206;
  rom[29738] = 16'hf1e6;
  rom[29739] = 16'hf227;
  rom[29740] = 16'hea07;
  rom[29741] = 16'hea28;
  rom[29742] = 16'hda48;
  rom[29743] = 16'hd247;
  rom[29744] = 16'hcac8;
  rom[29745] = 16'hc32a;
  rom[29746] = 16'hc34c;
  rom[29747] = 16'hcbcf;
  rom[29748] = 16'hd491;
  rom[29749] = 16'he533;
  rom[29750] = 16'hdd73;
  rom[29751] = 16'h82e6;
  rom[29752] = 16'hc54b;
  rom[29753] = 16'hf72f;
  rom[29754] = 16'hf70b;
  rom[29755] = 16'hff2a;
  rom[29756] = 16'hf709;
  rom[29757] = 16'hff2a;
  rom[29758] = 16'hef0c;
  rom[29759] = 16'hf70d;
  rom[29760] = 16'hef2d;
  rom[29761] = 16'hd66c;
  rom[29762] = 16'h5ac1;
  rom[29763] = 16'h8c0a;
  rom[29764] = 16'hf7bc;
  rom[29765] = 16'hffdf;
  rom[29766] = 16'hffbf;
  rom[29767] = 16'hffdf;
  rom[29768] = 16'hffff;
  rom[29769] = 16'hffff;
  rom[29770] = 16'hffff;
  rom[29771] = 16'hffff;
  rom[29772] = 16'hffff;
  rom[29773] = 16'hffff;
  rom[29774] = 16'hffff;
  rom[29775] = 16'hffff;
  rom[29776] = 16'hffff;
  rom[29777] = 16'hffff;
  rom[29778] = 16'hffff;
  rom[29779] = 16'hffff;
  rom[29780] = 16'hffff;
  rom[29781] = 16'hffff;
  rom[29782] = 16'hffff;
  rom[29783] = 16'hffff;
  rom[29784] = 16'hffff;
  rom[29785] = 16'hffff;
  rom[29786] = 16'hffff;
  rom[29787] = 16'hffff;
  rom[29788] = 16'hffff;
  rom[29789] = 16'hffff;
  rom[29790] = 16'hffff;
  rom[29791] = 16'hffff;
  rom[29792] = 16'hffff;
  rom[29793] = 16'hffff;
  rom[29794] = 16'hffff;
  rom[29795] = 16'hffff;
  rom[29796] = 16'hffff;
  rom[29797] = 16'hffff;
  rom[29798] = 16'hffff;
  rom[29799] = 16'hffff;
  rom[29800] = 16'hffff;
  rom[29801] = 16'hffff;
  rom[29802] = 16'hffff;
  rom[29803] = 16'hffff;
  rom[29804] = 16'hffff;
  rom[29805] = 16'hffff;
  rom[29806] = 16'hffff;
  rom[29807] = 16'hffff;
  rom[29808] = 16'hffff;
  rom[29809] = 16'hffff;
  rom[29810] = 16'hffff;
  rom[29811] = 16'hffff;
  rom[29812] = 16'hffff;
  rom[29813] = 16'hff1a;
  rom[29814] = 16'he450;
  rom[29815] = 16'hca47;
  rom[29816] = 16'hf248;
  rom[29817] = 16'he9c6;
  rom[29818] = 16'hfa27;
  rom[29819] = 16'hea26;
  rom[29820] = 16'hea27;
  rom[29821] = 16'hea26;
  rom[29822] = 16'hf227;
  rom[29823] = 16'hf207;
  rom[29824] = 16'hf227;
  rom[29825] = 16'hea07;
  rom[29826] = 16'hf228;
  rom[29827] = 16'hea06;
  rom[29828] = 16'hea26;
  rom[29829] = 16'hea26;
  rom[29830] = 16'hf227;
  rom[29831] = 16'hea06;
  rom[29832] = 16'hf226;
  rom[29833] = 16'hf206;
  rom[29834] = 16'hf247;
  rom[29835] = 16'hf206;
  rom[29836] = 16'hfa07;
  rom[29837] = 16'he207;
  rom[29838] = 16'hca88;
  rom[29839] = 16'h9243;
  rom[29840] = 16'hf66d;
  rom[29841] = 16'hfeea;
  rom[29842] = 16'hff29;
  rom[29843] = 16'hff08;
  rom[29844] = 16'hff2b;
  rom[29845] = 16'hef0b;
  rom[29846] = 16'hf72c;
  rom[29847] = 16'hf6cc;
  rom[29848] = 16'hc4a7;
  rom[29849] = 16'h81e1;
  rom[29850] = 16'hba66;
  rom[29851] = 16'hda69;
  rom[29852] = 16'hea48;
  rom[29853] = 16'he206;
  rom[29854] = 16'hf226;
  rom[29855] = 16'he9e5;
  rom[29856] = 16'hf227;
  rom[29857] = 16'hea07;
  rom[29858] = 16'hfa27;
  rom[29859] = 16'he9c5;
  rom[29860] = 16'hf247;
  rom[29861] = 16'he227;
  rom[29862] = 16'hd209;
  rom[29863] = 16'hc268;
  rom[29864] = 16'h91a4;
  rom[29865] = 16'h8aa2;
  rom[29866] = 16'hddcd;
  rom[29867] = 16'hd5ef;
  rom[29868] = 16'h7225;
  rom[29869] = 16'h89e6;
  rom[29870] = 16'hc2aa;
  rom[29871] = 16'hca88;
  rom[29872] = 16'hba46;
  rom[29873] = 16'ha1c3;
  rom[29874] = 16'h8963;
  rom[29875] = 16'h79a1;
  rom[29876] = 16'h8a84;
  rom[29877] = 16'ha407;
  rom[29878] = 16'hc4c9;
  rom[29879] = 16'he56b;
  rom[29880] = 16'hfe6e;
  rom[29881] = 16'hfe8b;
  rom[29882] = 16'hfeec;
  rom[29883] = 16'hf72d;
  rom[29884] = 16'hee4c;
  rom[29885] = 16'h92c3;
  rom[29886] = 16'ha9e3;
  rom[29887] = 16'hd267;
  rom[29888] = 16'hda87;
  rom[29889] = 16'hdaa7;
  rom[29890] = 16'hfcac;
  rom[29891] = 16'hec28;
  rom[29892] = 16'hf488;
  rom[29893] = 16'hd384;
  rom[29894] = 16'hcaa3;
  rom[29895] = 16'hdae6;
  rom[29896] = 16'hda86;
  rom[29897] = 16'hd285;
  rom[29898] = 16'hcac5;
  rom[29899] = 16'hbaa2;
  rom[29900] = 16'hdbc6;
  rom[29901] = 16'hec89;
  rom[29902] = 16'hf4cb;
  rom[29903] = 16'hf3c8;
  rom[29904] = 16'hdac6;
  rom[29905] = 16'hca65;
  rom[29906] = 16'hcaa6;
  rom[29907] = 16'h99e2;
  rom[29908] = 16'hab45;
  rom[29909] = 16'hf66b;
  rom[29910] = 16'hff6c;
  rom[29911] = 16'hf72a;
  rom[29912] = 16'hef2a;
  rom[29913] = 16'hef0b;
  rom[29914] = 16'hf70d;
  rom[29915] = 16'hf6ed;
  rom[29916] = 16'he66d;
  rom[29917] = 16'hcdca;
  rom[29918] = 16'hbd28;
  rom[29919] = 16'ha4a5;
  rom[29920] = 16'hc589;
  rom[29921] = 16'hd60b;
  rom[29922] = 16'hf6ef;
  rom[29923] = 16'hfeef;
  rom[29924] = 16'hcd4b;
  rom[29925] = 16'h79c0;
  rom[29926] = 16'hba66;
  rom[29927] = 16'hea47;
  rom[29928] = 16'hf1e6;
  rom[29929] = 16'hf205;
  rom[29930] = 16'hf227;
  rom[29931] = 16'he9e7;
  rom[29932] = 16'hf228;
  rom[29933] = 16'hf207;
  rom[29934] = 16'hf207;
  rom[29935] = 16'hf227;
  rom[29936] = 16'hea26;
  rom[29937] = 16'he206;
  rom[29938] = 16'hea28;
  rom[29939] = 16'he248;
  rom[29940] = 16'hda69;
  rom[29941] = 16'hd2ea;
  rom[29942] = 16'hdbee;
  rom[29943] = 16'hdcd1;
  rom[29944] = 16'hf5d5;
  rom[29945] = 16'hf678;
  rom[29946] = 16'hff3c;
  rom[29947] = 16'hff7d;
  rom[29948] = 16'hff5e;
  rom[29949] = 16'hff7d;
  rom[29950] = 16'hffbd;
  rom[29951] = 16'ha42c;
  rom[29952] = 16'h8386;
  rom[29953] = 16'hde6e;
  rom[29954] = 16'hf70e;
  rom[29955] = 16'hef2d;
  rom[29956] = 16'hf74d;
  rom[29957] = 16'hef2d;
  rom[29958] = 16'hf72f;
  rom[29959] = 16'he6cf;
  rom[29960] = 16'had0a;
  rom[29961] = 16'h5aa3;
  rom[29962] = 16'h944c;
  rom[29963] = 16'hef5a;
  rom[29964] = 16'hffff;
  rom[29965] = 16'hffff;
  rom[29966] = 16'hffff;
  rom[29967] = 16'hffff;
  rom[29968] = 16'hffff;
  rom[29969] = 16'hffff;
  rom[29970] = 16'hffff;
  rom[29971] = 16'hffff;
  rom[29972] = 16'hffff;
  rom[29973] = 16'hffff;
  rom[29974] = 16'hffff;
  rom[29975] = 16'hffff;
  rom[29976] = 16'hffff;
  rom[29977] = 16'hffff;
  rom[29978] = 16'hffff;
  rom[29979] = 16'hffff;
  rom[29980] = 16'hffff;
  rom[29981] = 16'hffff;
  rom[29982] = 16'hffff;
  rom[29983] = 16'hffff;
  rom[29984] = 16'hffff;
  rom[29985] = 16'hffff;
  rom[29986] = 16'hffff;
  rom[29987] = 16'hffff;
  rom[29988] = 16'hffff;
  rom[29989] = 16'hffff;
  rom[29990] = 16'hffff;
  rom[29991] = 16'hffff;
  rom[29992] = 16'hffff;
  rom[29993] = 16'hffff;
  rom[29994] = 16'hffff;
  rom[29995] = 16'hffff;
  rom[29996] = 16'hffff;
  rom[29997] = 16'hffff;
  rom[29998] = 16'hffff;
  rom[29999] = 16'hffff;
  rom[30000] = 16'hffff;
  rom[30001] = 16'hffff;
  rom[30002] = 16'hffff;
  rom[30003] = 16'hffff;
  rom[30004] = 16'hffff;
  rom[30005] = 16'hffff;
  rom[30006] = 16'hffff;
  rom[30007] = 16'hffff;
  rom[30008] = 16'hffff;
  rom[30009] = 16'hffff;
  rom[30010] = 16'hffff;
  rom[30011] = 16'hffff;
  rom[30012] = 16'hffde;
  rom[30013] = 16'hffde;
  rom[30014] = 16'hfe16;
  rom[30015] = 16'hd34c;
  rom[30016] = 16'hda28;
  rom[30017] = 16'hfa68;
  rom[30018] = 16'he1e5;
  rom[30019] = 16'hea26;
  rom[30020] = 16'hea46;
  rom[30021] = 16'he226;
  rom[30022] = 16'hea27;
  rom[30023] = 16'hf207;
  rom[30024] = 16'hf207;
  rom[30025] = 16'hf207;
  rom[30026] = 16'hea07;
  rom[30027] = 16'hea26;
  rom[30028] = 16'hea26;
  rom[30029] = 16'hea26;
  rom[30030] = 16'he226;
  rom[30031] = 16'hea06;
  rom[30032] = 16'hea06;
  rom[30033] = 16'hea26;
  rom[30034] = 16'he205;
  rom[30035] = 16'hf1e5;
  rom[30036] = 16'hf207;
  rom[30037] = 16'he228;
  rom[30038] = 16'hc287;
  rom[30039] = 16'h8a02;
  rom[30040] = 16'hee4d;
  rom[30041] = 16'hff0b;
  rom[30042] = 16'hff49;
  rom[30043] = 16'hff69;
  rom[30044] = 16'hf708;
  rom[30045] = 16'hef09;
  rom[30046] = 16'hef29;
  rom[30047] = 16'hff8c;
  rom[30048] = 16'hff2e;
  rom[30049] = 16'ha346;
  rom[30050] = 16'h89e2;
  rom[30051] = 16'hd289;
  rom[30052] = 16'hda27;
  rom[30053] = 16'hf268;
  rom[30054] = 16'hf246;
  rom[30055] = 16'hfa27;
  rom[30056] = 16'hf207;
  rom[30057] = 16'he9c7;
  rom[30058] = 16'he9c6;
  rom[30059] = 16'hfaa9;
  rom[30060] = 16'hd9e5;
  rom[30061] = 16'hda68;
  rom[30062] = 16'hc2a8;
  rom[30063] = 16'h91c3;
  rom[30064] = 16'h8a41;
  rom[30065] = 16'hd56a;
  rom[30066] = 16'hf70e;
  rom[30067] = 16'he68e;
  rom[30068] = 16'h72c6;
  rom[30069] = 16'h71c3;
  rom[30070] = 16'h81a2;
  rom[30071] = 16'h7920;
  rom[30072] = 16'h7920;
  rom[30073] = 16'ha2e4;
  rom[30074] = 16'he50b;
  rom[30075] = 16'hfeb0;
  rom[30076] = 16'hf6ae;
  rom[30077] = 16'hff2e;
  rom[30078] = 16'heeab;
  rom[30079] = 16'hf6cb;
  rom[30080] = 16'hfeea;
  rom[30081] = 16'hff4a;
  rom[30082] = 16'hf728;
  rom[30083] = 16'hf729;
  rom[30084] = 16'hf70c;
  rom[30085] = 16'hcd29;
  rom[30086] = 16'h7960;
  rom[30087] = 16'hba86;
  rom[30088] = 16'hd288;
  rom[30089] = 16'hd246;
  rom[30090] = 16'hdb06;
  rom[30091] = 16'hfd0d;
  rom[30092] = 16'he3a7;
  rom[30093] = 16'hc2a5;
  rom[30094] = 16'hdb07;
  rom[30095] = 16'hda87;
  rom[30096] = 16'heac8;
  rom[30097] = 16'heb08;
  rom[30098] = 16'hd2a6;
  rom[30099] = 16'he367;
  rom[30100] = 16'hd346;
  rom[30101] = 16'hec2a;
  rom[30102] = 16'hfc6b;
  rom[30103] = 16'hdac6;
  rom[30104] = 16'hca44;
  rom[30105] = 16'hca85;
  rom[30106] = 16'h9a43;
  rom[30107] = 16'h79c0;
  rom[30108] = 16'hddaa;
  rom[30109] = 16'hff4d;
  rom[30110] = 16'he6c9;
  rom[30111] = 16'hf72b;
  rom[30112] = 16'hff8e;
  rom[30113] = 16'hf70d;
  rom[30114] = 16'hc5a9;
  rom[30115] = 16'h7b62;
  rom[30116] = 16'h3960;
  rom[30117] = 16'h62a1;
  rom[30118] = 16'h9c45;
  rom[30119] = 16'hbd48;
  rom[30120] = 16'h83c3;
  rom[30121] = 16'h49e0;
  rom[30122] = 16'h6ac2;
  rom[30123] = 16'hcdcd;
  rom[30124] = 16'h9bc5;
  rom[30125] = 16'h9223;
  rom[30126] = 16'hc266;
  rom[30127] = 16'hea27;
  rom[30128] = 16'hf206;
  rom[30129] = 16'hf226;
  rom[30130] = 16'he206;
  rom[30131] = 16'hf227;
  rom[30132] = 16'hfa07;
  rom[30133] = 16'hf1c6;
  rom[30134] = 16'he9e7;
  rom[30135] = 16'he248;
  rom[30136] = 16'hda68;
  rom[30137] = 16'hda89;
  rom[30138] = 16'hca89;
  rom[30139] = 16'hdb6c;
  rom[30140] = 16'hf513;
  rom[30141] = 16'hfe98;
  rom[30142] = 16'hff7b;
  rom[30143] = 16'hffbd;
  rom[30144] = 16'hffde;
  rom[30145] = 16'hffde;
  rom[30146] = 16'hffbe;
  rom[30147] = 16'hffff;
  rom[30148] = 16'hffff;
  rom[30149] = 16'hffbf;
  rom[30150] = 16'hffbe;
  rom[30151] = 16'he6d9;
  rom[30152] = 16'h4203;
  rom[30153] = 16'h62e3;
  rom[30154] = 16'hb56b;
  rom[30155] = 16'hdecf;
  rom[30156] = 16'hc64d;
  rom[30157] = 16'hce2e;
  rom[30158] = 16'h9447;
  rom[30159] = 16'h4a01;
  rom[30160] = 16'h49e1;
  rom[30161] = 16'hbd71;
  rom[30162] = 16'hffbd;
  rom[30163] = 16'hffff;
  rom[30164] = 16'hffff;
  rom[30165] = 16'hffff;
  rom[30166] = 16'hffff;
  rom[30167] = 16'hffff;
  rom[30168] = 16'hffff;
  rom[30169] = 16'hffff;
  rom[30170] = 16'hffff;
  rom[30171] = 16'hffff;
  rom[30172] = 16'hffff;
  rom[30173] = 16'hffff;
  rom[30174] = 16'hffff;
  rom[30175] = 16'hffff;
  rom[30176] = 16'hffff;
  rom[30177] = 16'hffff;
  rom[30178] = 16'hffff;
  rom[30179] = 16'hffff;
  rom[30180] = 16'hffff;
  rom[30181] = 16'hffff;
  rom[30182] = 16'hffff;
  rom[30183] = 16'hffff;
  rom[30184] = 16'hffff;
  rom[30185] = 16'hffff;
  rom[30186] = 16'hffff;
  rom[30187] = 16'hffff;
  rom[30188] = 16'hffff;
  rom[30189] = 16'hffff;
  rom[30190] = 16'hffff;
  rom[30191] = 16'hffff;
  rom[30192] = 16'hffff;
  rom[30193] = 16'hffff;
  rom[30194] = 16'hffff;
  rom[30195] = 16'hffff;
  rom[30196] = 16'hffff;
  rom[30197] = 16'hffff;
  rom[30198] = 16'hffff;
  rom[30199] = 16'hffff;
  rom[30200] = 16'hffff;
  rom[30201] = 16'hffff;
  rom[30202] = 16'hffff;
  rom[30203] = 16'hffff;
  rom[30204] = 16'hffff;
  rom[30205] = 16'hffff;
  rom[30206] = 16'hffff;
  rom[30207] = 16'hffff;
  rom[30208] = 16'hffff;
  rom[30209] = 16'hffff;
  rom[30210] = 16'hffff;
  rom[30211] = 16'hffff;
  rom[30212] = 16'hffff;
  rom[30213] = 16'hffdf;
  rom[30214] = 16'hff1c;
  rom[30215] = 16'hecb1;
  rom[30216] = 16'hd269;
  rom[30217] = 16'he227;
  rom[30218] = 16'hea26;
  rom[30219] = 16'hea46;
  rom[30220] = 16'hea46;
  rom[30221] = 16'he246;
  rom[30222] = 16'hea27;
  rom[30223] = 16'hf207;
  rom[30224] = 16'hf228;
  rom[30225] = 16'hf207;
  rom[30226] = 16'hf227;
  rom[30227] = 16'hea06;
  rom[30228] = 16'hea47;
  rom[30229] = 16'hea26;
  rom[30230] = 16'hea46;
  rom[30231] = 16'hea06;
  rom[30232] = 16'hf227;
  rom[30233] = 16'hea26;
  rom[30234] = 16'hf246;
  rom[30235] = 16'hea06;
  rom[30236] = 16'hfa47;
  rom[30237] = 16'he207;
  rom[30238] = 16'hd267;
  rom[30239] = 16'h89c2;
  rom[30240] = 16'he58c;
  rom[30241] = 16'hfeec;
  rom[30242] = 16'hf729;
  rom[30243] = 16'heee7;
  rom[30244] = 16'hff69;
  rom[30245] = 16'hf728;
  rom[30246] = 16'hff4a;
  rom[30247] = 16'hef29;
  rom[30248] = 16'hff0c;
  rom[30249] = 16'hee2c;
  rom[30250] = 16'h8a42;
  rom[30251] = 16'h99c3;
  rom[30252] = 16'hd268;
  rom[30253] = 16'he228;
  rom[30254] = 16'hea07;
  rom[30255] = 16'hf247;
  rom[30256] = 16'hf229;
  rom[30257] = 16'hea29;
  rom[30258] = 16'hea29;
  rom[30259] = 16'hd1e6;
  rom[30260] = 16'hd287;
  rom[30261] = 16'hb224;
  rom[30262] = 16'h91c1;
  rom[30263] = 16'h92a3;
  rom[30264] = 16'hfe6d;
  rom[30265] = 16'hfeec;
  rom[30266] = 16'hff0b;
  rom[30267] = 16'heecc;
  rom[30268] = 16'h8be6;
  rom[30269] = 16'h51c0;
  rom[30270] = 16'ha3e6;
  rom[30271] = 16'hcd09;
  rom[30272] = 16'hfeae;
  rom[30273] = 16'hfead;
  rom[30274] = 16'hfeed;
  rom[30275] = 16'hfecc;
  rom[30276] = 16'hff0b;
  rom[30277] = 16'hff0a;
  rom[30278] = 16'hff29;
  rom[30279] = 16'hff0a;
  rom[30280] = 16'hff2a;
  rom[30281] = 16'hff07;
  rom[30282] = 16'hff28;
  rom[30283] = 16'hf707;
  rom[30284] = 16'hff4c;
  rom[30285] = 16'hf6ad;
  rom[30286] = 16'hc489;
  rom[30287] = 16'h8a02;
  rom[30288] = 16'hba86;
  rom[30289] = 16'hcaa6;
  rom[30290] = 16'hd2c6;
  rom[30291] = 16'hebca;
  rom[30292] = 16'hf42c;
  rom[30293] = 16'hfc0c;
  rom[30294] = 16'hfc0c;
  rom[30295] = 16'hf3cb;
  rom[30296] = 16'hfc0c;
  rom[30297] = 16'hfbeb;
  rom[30298] = 16'hfc2c;
  rom[30299] = 16'hf3ea;
  rom[30300] = 16'hfc0a;
  rom[30301] = 16'hf42c;
  rom[30302] = 16'hf3aa;
  rom[30303] = 16'hd2a6;
  rom[30304] = 16'hd2c6;
  rom[30305] = 16'hb284;
  rom[30306] = 16'h8a01;
  rom[30307] = 16'hcce8;
  rom[30308] = 16'hfeee;
  rom[30309] = 16'hf70d;
  rom[30310] = 16'hef0d;
  rom[30311] = 16'he6ac;
  rom[30312] = 16'hb506;
  rom[30313] = 16'h83c2;
  rom[30314] = 16'h83a5;
  rom[30315] = 16'hb548;
  rom[30316] = 16'hf6cf;
  rom[30317] = 16'heeee;
  rom[30318] = 16'hef0d;
  rom[30319] = 16'hef0c;
  rom[30320] = 16'hef0d;
  rom[30321] = 16'hef0f;
  rom[30322] = 16'hace9;
  rom[30323] = 16'h8345;
  rom[30324] = 16'h7224;
  rom[30325] = 16'h89e4;
  rom[30326] = 16'hd269;
  rom[30327] = 16'hea08;
  rom[30328] = 16'hf208;
  rom[30329] = 16'hea26;
  rom[30330] = 16'hea47;
  rom[30331] = 16'hf227;
  rom[30332] = 16'hf9e7;
  rom[30333] = 16'hf207;
  rom[30334] = 16'hea49;
  rom[30335] = 16'hd268;
  rom[30336] = 16'hd2ea;
  rom[30337] = 16'hdbee;
  rom[30338] = 16'hf575;
  rom[30339] = 16'hfeb9;
  rom[30340] = 16'hff7d;
  rom[30341] = 16'hffdd;
  rom[30342] = 16'hffff;
  rom[30343] = 16'hffff;
  rom[30344] = 16'hffff;
  rom[30345] = 16'hffdf;
  rom[30346] = 16'hffdf;
  rom[30347] = 16'hffdf;
  rom[30348] = 16'hffdf;
  rom[30349] = 16'hffdf;
  rom[30350] = 16'hffff;
  rom[30351] = 16'hffde;
  rom[30352] = 16'hd677;
  rom[30353] = 16'h9cce;
  rom[30354] = 16'h7bc9;
  rom[30355] = 16'h6305;
  rom[30356] = 16'h6306;
  rom[30357] = 16'h6b47;
  rom[30358] = 16'h8c0b;
  rom[30359] = 16'had10;
  rom[30360] = 16'he6d9;
  rom[30361] = 16'hffde;
  rom[30362] = 16'hffff;
  rom[30363] = 16'hffff;
  rom[30364] = 16'hffff;
  rom[30365] = 16'hffff;
  rom[30366] = 16'hffff;
  rom[30367] = 16'hffff;
  rom[30368] = 16'hffff;
  rom[30369] = 16'hffff;
  rom[30370] = 16'hffff;
  rom[30371] = 16'hffff;
  rom[30372] = 16'hffff;
  rom[30373] = 16'hffff;
  rom[30374] = 16'hffff;
  rom[30375] = 16'hffff;
  rom[30376] = 16'hffff;
  rom[30377] = 16'hffff;
  rom[30378] = 16'hffff;
  rom[30379] = 16'hffff;
  rom[30380] = 16'hffff;
  rom[30381] = 16'hffff;
  rom[30382] = 16'hffff;
  rom[30383] = 16'hffff;
  rom[30384] = 16'hffff;
  rom[30385] = 16'hffff;
  rom[30386] = 16'hffff;
  rom[30387] = 16'hffff;
  rom[30388] = 16'hffff;
  rom[30389] = 16'hffff;
  rom[30390] = 16'hffff;
  rom[30391] = 16'hffff;
  rom[30392] = 16'hffff;
  rom[30393] = 16'hffff;
  rom[30394] = 16'hffff;
  rom[30395] = 16'hffff;
  rom[30396] = 16'hffff;
  rom[30397] = 16'hffff;
  rom[30398] = 16'hffff;
  rom[30399] = 16'hffff;
  rom[30400] = 16'hffff;
  rom[30401] = 16'hffff;
  rom[30402] = 16'hffff;
  rom[30403] = 16'hffff;
  rom[30404] = 16'hffff;
  rom[30405] = 16'hffff;
  rom[30406] = 16'hffff;
  rom[30407] = 16'hffff;
  rom[30408] = 16'hffff;
  rom[30409] = 16'hffff;
  rom[30410] = 16'hffff;
  rom[30411] = 16'hffff;
  rom[30412] = 16'hffdf;
  rom[30413] = 16'hffff;
  rom[30414] = 16'hff9e;
  rom[30415] = 16'hfeb9;
  rom[30416] = 16'hd3ac;
  rom[30417] = 16'hd246;
  rom[30418] = 16'hea66;
  rom[30419] = 16'hea45;
  rom[30420] = 16'hea25;
  rom[30421] = 16'hea46;
  rom[30422] = 16'hea26;
  rom[30423] = 16'hf1e7;
  rom[30424] = 16'hea07;
  rom[30425] = 16'hf207;
  rom[30426] = 16'hf227;
  rom[30427] = 16'hea26;
  rom[30428] = 16'he226;
  rom[30429] = 16'hea26;
  rom[30430] = 16'hea26;
  rom[30431] = 16'hea06;
  rom[30432] = 16'hea06;
  rom[30433] = 16'hea06;
  rom[30434] = 16'hea26;
  rom[30435] = 16'hea26;
  rom[30436] = 16'hea26;
  rom[30437] = 16'hea26;
  rom[30438] = 16'hd267;
  rom[30439] = 16'ha1e3;
  rom[30440] = 16'hb3e7;
  rom[30441] = 16'hf70e;
  rom[30442] = 16'hef4b;
  rom[30443] = 16'he728;
  rom[30444] = 16'hf748;
  rom[30445] = 16'hff08;
  rom[30446] = 16'hff08;
  rom[30447] = 16'hf708;
  rom[30448] = 16'hef2a;
  rom[30449] = 16'hff0c;
  rom[30450] = 16'he5cb;
  rom[30451] = 16'h9201;
  rom[30452] = 16'hb225;
  rom[30453] = 16'hca47;
  rom[30454] = 16'hda88;
  rom[30455] = 16'hda47;
  rom[30456] = 16'hda47;
  rom[30457] = 16'hda68;
  rom[30458] = 16'hca67;
  rom[30459] = 16'hd2c8;
  rom[30460] = 16'h99e2;
  rom[30461] = 16'h89a0;
  rom[30462] = 16'hbc26;
  rom[30463] = 16'hfe6c;
  rom[30464] = 16'hfeca;
  rom[30465] = 16'hf6c9;
  rom[30466] = 16'hf6c9;
  rom[30467] = 16'hfeed;
  rom[30468] = 16'hb54a;
  rom[30469] = 16'h5200;
  rom[30470] = 16'hc5aa;
  rom[30471] = 16'heecc;
  rom[30472] = 16'hff2a;
  rom[30473] = 16'hff4b;
  rom[30474] = 16'hff0a;
  rom[30475] = 16'hff0a;
  rom[30476] = 16'hff29;
  rom[30477] = 16'hff49;
  rom[30478] = 16'hff08;
  rom[30479] = 16'hff29;
  rom[30480] = 16'hff08;
  rom[30481] = 16'hff07;
  rom[30482] = 16'hff07;
  rom[30483] = 16'hfee7;
  rom[30484] = 16'hf6ea;
  rom[30485] = 16'hf6ed;
  rom[30486] = 16'hf6ce;
  rom[30487] = 16'hbc48;
  rom[30488] = 16'h79c0;
  rom[30489] = 16'ha222;
  rom[30490] = 16'hc265;
  rom[30491] = 16'hdaa7;
  rom[30492] = 16'hdaa7;
  rom[30493] = 16'hdaa7;
  rom[30494] = 16'hda66;
  rom[30495] = 16'he287;
  rom[30496] = 16'hda65;
  rom[30497] = 16'he265;
  rom[30498] = 16'he2a6;
  rom[30499] = 16'hda66;
  rom[30500] = 16'he2a7;
  rom[30501] = 16'hdac8;
  rom[30502] = 16'hcaa8;
  rom[30503] = 16'hcaa6;
  rom[30504] = 16'h91a1;
  rom[30505] = 16'h9221;
  rom[30506] = 16'hc468;
  rom[30507] = 16'hff0f;
  rom[30508] = 16'heeed;
  rom[30509] = 16'hef0e;
  rom[30510] = 16'hc5c9;
  rom[30511] = 16'h8bc3;
  rom[30512] = 16'h83a0;
  rom[30513] = 16'hcde8;
  rom[30514] = 16'hef0c;
  rom[30515] = 16'hf70d;
  rom[30516] = 16'hf70c;
  rom[30517] = 16'hf72a;
  rom[30518] = 16'hef08;
  rom[30519] = 16'hf728;
  rom[30520] = 16'hf729;
  rom[30521] = 16'hff6d;
  rom[30522] = 16'heeee;
  rom[30523] = 16'hd5cd;
  rom[30524] = 16'h8b05;
  rom[30525] = 16'h89c4;
  rom[30526] = 16'hd28a;
  rom[30527] = 16'he208;
  rom[30528] = 16'hea48;
  rom[30529] = 16'hea27;
  rom[30530] = 16'he227;
  rom[30531] = 16'hf206;
  rom[30532] = 16'he9c5;
  rom[30533] = 16'hf289;
  rom[30534] = 16'hca68;
  rom[30535] = 16'hd36d;
  rom[30536] = 16'hf554;
  rom[30537] = 16'hfefb;
  rom[30538] = 16'hff7c;
  rom[30539] = 16'hfffe;
  rom[30540] = 16'hffde;
  rom[30541] = 16'hffff;
  rom[30542] = 16'hffbe;
  rom[30543] = 16'hffff;
  rom[30544] = 16'hffdf;
  rom[30545] = 16'hffdf;
  rom[30546] = 16'hffdf;
  rom[30547] = 16'hffff;
  rom[30548] = 16'hffdf;
  rom[30549] = 16'hffff;
  rom[30550] = 16'hffdf;
  rom[30551] = 16'hffff;
  rom[30552] = 16'hfffe;
  rom[30553] = 16'hfffe;
  rom[30554] = 16'hf7bc;
  rom[30555] = 16'hf77b;
  rom[30556] = 16'hef5b;
  rom[30557] = 16'hf75b;
  rom[30558] = 16'hffdd;
  rom[30559] = 16'hffff;
  rom[30560] = 16'hffdf;
  rom[30561] = 16'hffdf;
  rom[30562] = 16'hffdf;
  rom[30563] = 16'hffff;
  rom[30564] = 16'hffff;
  rom[30565] = 16'hffff;
  rom[30566] = 16'hffff;
  rom[30567] = 16'hffff;
  rom[30568] = 16'hffff;
  rom[30569] = 16'hffff;
  rom[30570] = 16'hffff;
  rom[30571] = 16'hffff;
  rom[30572] = 16'hffff;
  rom[30573] = 16'hffff;
  rom[30574] = 16'hffff;
  rom[30575] = 16'hffff;
  rom[30576] = 16'hffff;
  rom[30577] = 16'hffff;
  rom[30578] = 16'hffff;
  rom[30579] = 16'hffff;
  rom[30580] = 16'hffff;
  rom[30581] = 16'hffff;
  rom[30582] = 16'hffff;
  rom[30583] = 16'hffff;
  rom[30584] = 16'hffff;
  rom[30585] = 16'hffff;
  rom[30586] = 16'hffff;
  rom[30587] = 16'hffff;
  rom[30588] = 16'hffff;
  rom[30589] = 16'hffff;
  rom[30590] = 16'hffff;
  rom[30591] = 16'hffff;
  rom[30592] = 16'hffff;
  rom[30593] = 16'hffff;
  rom[30594] = 16'hffff;
  rom[30595] = 16'hffff;
  rom[30596] = 16'hffff;
  rom[30597] = 16'hffff;
  rom[30598] = 16'hffff;
  rom[30599] = 16'hffff;
  rom[30600] = 16'hffff;
  rom[30601] = 16'hffff;
  rom[30602] = 16'hffff;
  rom[30603] = 16'hffff;
  rom[30604] = 16'hffff;
  rom[30605] = 16'hffff;
  rom[30606] = 16'hffff;
  rom[30607] = 16'hffff;
  rom[30608] = 16'hffff;
  rom[30609] = 16'hffff;
  rom[30610] = 16'hffff;
  rom[30611] = 16'hffff;
  rom[30612] = 16'hffff;
  rom[30613] = 16'hffff;
  rom[30614] = 16'hffff;
  rom[30615] = 16'hff9d;
  rom[30616] = 16'hfdd6;
  rom[30617] = 16'hc329;
  rom[30618] = 16'hda67;
  rom[30619] = 16'hea46;
  rom[30620] = 16'hf226;
  rom[30621] = 16'hf206;
  rom[30622] = 16'hfa27;
  rom[30623] = 16'hf207;
  rom[30624] = 16'hf227;
  rom[30625] = 16'hf207;
  rom[30626] = 16'hf228;
  rom[30627] = 16'hea26;
  rom[30628] = 16'hea26;
  rom[30629] = 16'hea26;
  rom[30630] = 16'hea27;
  rom[30631] = 16'hea06;
  rom[30632] = 16'hf226;
  rom[30633] = 16'hea07;
  rom[30634] = 16'hf248;
  rom[30635] = 16'hea26;
  rom[30636] = 16'hf266;
  rom[30637] = 16'hea25;
  rom[30638] = 16'he288;
  rom[30639] = 16'hb204;
  rom[30640] = 16'h8a22;
  rom[30641] = 16'hde2d;
  rom[30642] = 16'hef4e;
  rom[30643] = 16'hef6a;
  rom[30644] = 16'hf768;
  rom[30645] = 16'hff28;
  rom[30646] = 16'hfee8;
  rom[30647] = 16'hff49;
  rom[30648] = 16'hf709;
  rom[30649] = 16'hef2a;
  rom[30650] = 16'hfeec;
  rom[30651] = 16'hd4e9;
  rom[30652] = 16'h8a21;
  rom[30653] = 16'h99e3;
  rom[30654] = 16'hba46;
  rom[30655] = 16'hc2a6;
  rom[30656] = 16'hc286;
  rom[30657] = 16'hbaa5;
  rom[30658] = 16'ha223;
  rom[30659] = 16'h89e0;
  rom[30660] = 16'h9ac3;
  rom[30661] = 16'hd508;
  rom[30662] = 16'hfecc;
  rom[30663] = 16'hfeea;
  rom[30664] = 16'hff29;
  rom[30665] = 16'hff4b;
  rom[30666] = 16'hff0c;
  rom[30667] = 16'hf6ee;
  rom[30668] = 16'haca9;
  rom[30669] = 16'h4180;
  rom[30670] = 16'hbd69;
  rom[30671] = 16'hff8e;
  rom[30672] = 16'hf709;
  rom[30673] = 16'hf708;
  rom[30674] = 16'hff2a;
  rom[30675] = 16'hff49;
  rom[30676] = 16'hff08;
  rom[30677] = 16'hf6e7;
  rom[30678] = 16'hff29;
  rom[30679] = 16'hf729;
  rom[30680] = 16'hff2a;
  rom[30681] = 16'hf708;
  rom[30682] = 16'hff29;
  rom[30683] = 16'hfee7;
  rom[30684] = 16'hff2a;
  rom[30685] = 16'hf70b;
  rom[30686] = 16'hff2d;
  rom[30687] = 16'hee8d;
  rom[30688] = 16'hbca7;
  rom[30689] = 16'h8a41;
  rom[30690] = 16'ha1c1;
  rom[30691] = 16'hca65;
  rom[30692] = 16'hd266;
  rom[30693] = 16'hd266;
  rom[30694] = 16'he287;
  rom[30695] = 16'hda66;
  rom[30696] = 16'hda66;
  rom[30697] = 16'hda46;
  rom[30698] = 16'he287;
  rom[30699] = 16'hda87;
  rom[30700] = 16'hd287;
  rom[30701] = 16'hc265;
  rom[30702] = 16'hb245;
  rom[30703] = 16'h9a23;
  rom[30704] = 16'h9aa3;
  rom[30705] = 16'hcce8;
  rom[30706] = 16'hfeef;
  rom[30707] = 16'hfeee;
  rom[30708] = 16'he6ad;
  rom[30709] = 16'had28;
  rom[30710] = 16'h83a3;
  rom[30711] = 16'hacc6;
  rom[30712] = 16'hff0d;
  rom[30713] = 16'hff4b;
  rom[30714] = 16'hf70a;
  rom[30715] = 16'hf70a;
  rom[30716] = 16'hf709;
  rom[30717] = 16'hf728;
  rom[30718] = 16'hff48;
  rom[30719] = 16'hff87;
  rom[30720] = 16'hf727;
  rom[30721] = 16'hf708;
  rom[30722] = 16'hf72c;
  rom[30723] = 16'hff0e;
  rom[30724] = 16'hd52b;
  rom[30725] = 16'h9a85;
  rom[30726] = 16'hc248;
  rom[30727] = 16'he249;
  rom[30728] = 16'he228;
  rom[30729] = 16'he226;
  rom[30730] = 16'hea27;
  rom[30731] = 16'he9e6;
  rom[30732] = 16'hf267;
  rom[30733] = 16'hd247;
  rom[30734] = 16'hd3ce;
  rom[30735] = 16'hfe17;
  rom[30736] = 16'hff7d;
  rom[30737] = 16'hffbe;
  rom[30738] = 16'hffdf;
  rom[30739] = 16'hffff;
  rom[30740] = 16'hffff;
  rom[30741] = 16'hffdf;
  rom[30742] = 16'hffbf;
  rom[30743] = 16'hffbf;
  rom[30744] = 16'hffff;
  rom[30745] = 16'hffff;
  rom[30746] = 16'hffff;
  rom[30747] = 16'hffff;
  rom[30748] = 16'hffdf;
  rom[30749] = 16'hffdf;
  rom[30750] = 16'hffdf;
  rom[30751] = 16'hffff;
  rom[30752] = 16'hffff;
  rom[30753] = 16'hffde;
  rom[30754] = 16'hffff;
  rom[30755] = 16'hffff;
  rom[30756] = 16'hffff;
  rom[30757] = 16'hffdf;
  rom[30758] = 16'hffdf;
  rom[30759] = 16'hffdf;
  rom[30760] = 16'hffdf;
  rom[30761] = 16'hffdf;
  rom[30762] = 16'hffff;
  rom[30763] = 16'hffff;
  rom[30764] = 16'hffff;
  rom[30765] = 16'hffff;
  rom[30766] = 16'hffff;
  rom[30767] = 16'hffff;
  rom[30768] = 16'hffff;
  rom[30769] = 16'hffff;
  rom[30770] = 16'hffff;
  rom[30771] = 16'hffff;
  rom[30772] = 16'hffff;
  rom[30773] = 16'hffff;
  rom[30774] = 16'hffff;
  rom[30775] = 16'hffff;
  rom[30776] = 16'hffff;
  rom[30777] = 16'hffff;
  rom[30778] = 16'hffff;
  rom[30779] = 16'hffff;
  rom[30780] = 16'hffff;
  rom[30781] = 16'hffff;
  rom[30782] = 16'hffff;
  rom[30783] = 16'hffff;
  rom[30784] = 16'hffff;
  rom[30785] = 16'hffff;
  rom[30786] = 16'hffff;
  rom[30787] = 16'hffff;
  rom[30788] = 16'hffff;
  rom[30789] = 16'hffff;
  rom[30790] = 16'hffff;
  rom[30791] = 16'hffff;
  rom[30792] = 16'hffff;
  rom[30793] = 16'hffff;
  rom[30794] = 16'hffff;
  rom[30795] = 16'hffff;
  rom[30796] = 16'hffff;
  rom[30797] = 16'hffff;
  rom[30798] = 16'hffff;
  rom[30799] = 16'hffff;
  rom[30800] = 16'hffff;
  rom[30801] = 16'hffff;
  rom[30802] = 16'hffff;
  rom[30803] = 16'hffff;
  rom[30804] = 16'hffff;
  rom[30805] = 16'hffff;
  rom[30806] = 16'hffff;
  rom[30807] = 16'hffff;
  rom[30808] = 16'hffff;
  rom[30809] = 16'hffff;
  rom[30810] = 16'hffff;
  rom[30811] = 16'hffff;
  rom[30812] = 16'hffff;
  rom[30813] = 16'hffff;
  rom[30814] = 16'hffff;
  rom[30815] = 16'hffdf;
  rom[30816] = 16'hff5b;
  rom[30817] = 16'hed32;
  rom[30818] = 16'hd329;
  rom[30819] = 16'hda26;
  rom[30820] = 16'he9e6;
  rom[30821] = 16'hf206;
  rom[30822] = 16'hf1e6;
  rom[30823] = 16'hf227;
  rom[30824] = 16'hea07;
  rom[30825] = 16'hf227;
  rom[30826] = 16'hea06;
  rom[30827] = 16'hf227;
  rom[30828] = 16'hea06;
  rom[30829] = 16'hea06;
  rom[30830] = 16'he206;
  rom[30831] = 16'hea06;
  rom[30832] = 16'hea06;
  rom[30833] = 16'hea07;
  rom[30834] = 16'hea07;
  rom[30835] = 16'hea26;
  rom[30836] = 16'hea46;
  rom[30837] = 16'hea45;
  rom[30838] = 16'he247;
  rom[30839] = 16'hca46;
  rom[30840] = 16'h8982;
  rom[30841] = 16'habe7;
  rom[30842] = 16'heeef;
  rom[30843] = 16'hdeca;
  rom[30844] = 16'hf74a;
  rom[30845] = 16'hf6c8;
  rom[30846] = 16'hff09;
  rom[30847] = 16'hff29;
  rom[30848] = 16'hf729;
  rom[30849] = 16'hf729;
  rom[30850] = 16'hef4a;
  rom[30851] = 16'hf6ec;
  rom[30852] = 16'he5cb;
  rom[30853] = 16'hb3c7;
  rom[30854] = 16'h8a41;
  rom[30855] = 16'h9241;
  rom[30856] = 16'h9280;
  rom[30857] = 16'h9280;
  rom[30858] = 16'ha382;
  rom[30859] = 16'hcce7;
  rom[30860] = 16'hee0b;
  rom[30861] = 16'hfecd;
  rom[30862] = 16'hf6e9;
  rom[30863] = 16'hff49;
  rom[30864] = 16'he6e8;
  rom[30865] = 16'hf74d;
  rom[30866] = 16'hef0e;
  rom[30867] = 16'hc50a;
  rom[30868] = 16'h7a42;
  rom[30869] = 16'h59c1;
  rom[30870] = 16'h9c26;
  rom[30871] = 16'hf72d;
  rom[30872] = 16'hf709;
  rom[30873] = 16'hff29;
  rom[30874] = 16'hf709;
  rom[30875] = 16'hff2a;
  rom[30876] = 16'hf729;
  rom[30877] = 16'hf729;
  rom[30878] = 16'hef09;
  rom[30879] = 16'hef4a;
  rom[30880] = 16'hef2a;
  rom[30881] = 16'hf72a;
  rom[30882] = 16'hff29;
  rom[30883] = 16'hff28;
  rom[30884] = 16'hf728;
  rom[30885] = 16'hff49;
  rom[30886] = 16'he709;
  rom[30887] = 16'hef0c;
  rom[30888] = 16'hf6ee;
  rom[30889] = 16'hdd8a;
  rom[30890] = 16'hbbc4;
  rom[30891] = 16'h9200;
  rom[30892] = 16'ha1c1;
  rom[30893] = 16'hb1e3;
  rom[30894] = 16'hba24;
  rom[30895] = 16'hca86;
  rom[30896] = 16'hc245;
  rom[30897] = 16'hc246;
  rom[30898] = 16'hba46;
  rom[30899] = 16'hb246;
  rom[30900] = 16'h99e2;
  rom[30901] = 16'h9a02;
  rom[30902] = 16'h9220;
  rom[30903] = 16'hb3c6;
  rom[30904] = 16'he60b;
  rom[30905] = 16'hff0d;
  rom[30906] = 16'hf6ec;
  rom[30907] = 16'heecd;
  rom[30908] = 16'h9c45;
  rom[30909] = 16'h83c4;
  rom[30910] = 16'hc5c9;
  rom[30911] = 16'heeed;
  rom[30912] = 16'hff0b;
  rom[30913] = 16'hff2a;
  rom[30914] = 16'hf729;
  rom[30915] = 16'hff29;
  rom[30916] = 16'hff29;
  rom[30917] = 16'hff29;
  rom[30918] = 16'hf707;
  rom[30919] = 16'hf707;
  rom[30920] = 16'hff48;
  rom[30921] = 16'hf708;
  rom[30922] = 16'hff2a;
  rom[30923] = 16'hff0c;
  rom[30924] = 16'hf66c;
  rom[30925] = 16'hb3a6;
  rom[30926] = 16'ha203;
  rom[30927] = 16'hd287;
  rom[30928] = 16'he226;
  rom[30929] = 16'hea26;
  rom[30930] = 16'he226;
  rom[30931] = 16'he226;
  rom[30932] = 16'hd247;
  rom[30933] = 16'hdb8c;
  rom[30934] = 16'hfe57;
  rom[30935] = 16'hff7d;
  rom[30936] = 16'hffde;
  rom[30937] = 16'hffff;
  rom[30938] = 16'hffff;
  rom[30939] = 16'hffff;
  rom[30940] = 16'hffff;
  rom[30941] = 16'hffff;
  rom[30942] = 16'hffff;
  rom[30943] = 16'hffff;
  rom[30944] = 16'hffff;
  rom[30945] = 16'hffff;
  rom[30946] = 16'hffff;
  rom[30947] = 16'hffff;
  rom[30948] = 16'hffff;
  rom[30949] = 16'hffff;
  rom[30950] = 16'hffff;
  rom[30951] = 16'hffff;
  rom[30952] = 16'hffff;
  rom[30953] = 16'hffff;
  rom[30954] = 16'hffff;
  rom[30955] = 16'hffff;
  rom[30956] = 16'hffff;
  rom[30957] = 16'hffff;
  rom[30958] = 16'hffff;
  rom[30959] = 16'hffff;
  rom[30960] = 16'hffdf;
  rom[30961] = 16'hffff;
  rom[30962] = 16'hffff;
  rom[30963] = 16'hffff;
  rom[30964] = 16'hffff;
  rom[30965] = 16'hffff;
  rom[30966] = 16'hffff;
  rom[30967] = 16'hffff;
  rom[30968] = 16'hffff;
  rom[30969] = 16'hffff;
  rom[30970] = 16'hffff;
  rom[30971] = 16'hffff;
  rom[30972] = 16'hffff;
  rom[30973] = 16'hffff;
  rom[30974] = 16'hffff;
  rom[30975] = 16'hffff;
  rom[30976] = 16'hffff;
  rom[30977] = 16'hffff;
  rom[30978] = 16'hffff;
  rom[30979] = 16'hffff;
  rom[30980] = 16'hffff;
  rom[30981] = 16'hffff;
  rom[30982] = 16'hffff;
  rom[30983] = 16'hffff;
  rom[30984] = 16'hffff;
  rom[30985] = 16'hffff;
  rom[30986] = 16'hffff;
  rom[30987] = 16'hffff;
  rom[30988] = 16'hffff;
  rom[30989] = 16'hffff;
  rom[30990] = 16'hffff;
  rom[30991] = 16'hffff;
  rom[30992] = 16'hffff;
  rom[30993] = 16'hffff;
  rom[30994] = 16'hffff;
  rom[30995] = 16'hffff;
  rom[30996] = 16'hffff;
  rom[30997] = 16'hffff;
  rom[30998] = 16'hffff;
  rom[30999] = 16'hffff;
  rom[31000] = 16'hffff;
  rom[31001] = 16'hffff;
  rom[31002] = 16'hffff;
  rom[31003] = 16'hffff;
  rom[31004] = 16'hffff;
  rom[31005] = 16'hffff;
  rom[31006] = 16'hffff;
  rom[31007] = 16'hffff;
  rom[31008] = 16'hffff;
  rom[31009] = 16'hffff;
  rom[31010] = 16'hffff;
  rom[31011] = 16'hffff;
  rom[31012] = 16'hffff;
  rom[31013] = 16'hffff;
  rom[31014] = 16'hffff;
  rom[31015] = 16'hfffe;
  rom[31016] = 16'hfffe;
  rom[31017] = 16'hfefa;
  rom[31018] = 16'he4d1;
  rom[31019] = 16'hdb0a;
  rom[31020] = 16'he248;
  rom[31021] = 16'he9e6;
  rom[31022] = 16'hf1e7;
  rom[31023] = 16'hea47;
  rom[31024] = 16'hea48;
  rom[31025] = 16'hea27;
  rom[31026] = 16'hea27;
  rom[31027] = 16'hf227;
  rom[31028] = 16'hf227;
  rom[31029] = 16'hf206;
  rom[31030] = 16'hf226;
  rom[31031] = 16'hea06;
  rom[31032] = 16'hea27;
  rom[31033] = 16'hea07;
  rom[31034] = 16'hea27;
  rom[31035] = 16'he206;
  rom[31036] = 16'hea67;
  rom[31037] = 16'he226;
  rom[31038] = 16'hea47;
  rom[31039] = 16'he247;
  rom[31040] = 16'hba26;
  rom[31041] = 16'h81e2;
  rom[31042] = 16'hd52b;
  rom[31043] = 16'hff8f;
  rom[31044] = 16'hf70b;
  rom[31045] = 16'hff4b;
  rom[31046] = 16'hf6c9;
  rom[31047] = 16'hff29;
  rom[31048] = 16'hf729;
  rom[31049] = 16'hf708;
  rom[31050] = 16'hf76a;
  rom[31051] = 16'hef0a;
  rom[31052] = 16'hf70d;
  rom[31053] = 16'hf6cd;
  rom[31054] = 16'hfece;
  rom[31055] = 16'hdd89;
  rom[31056] = 16'he5a9;
  rom[31057] = 16'hff0d;
  rom[31058] = 16'hfeca;
  rom[31059] = 16'hff2c;
  rom[31060] = 16'hff0c;
  rom[31061] = 16'hff2b;
  rom[31062] = 16'hf70a;
  rom[31063] = 16'hf76a;
  rom[31064] = 16'hf72b;
  rom[31065] = 16'hf70e;
  rom[31066] = 16'hd5ac;
  rom[31067] = 16'h7a01;
  rom[31068] = 16'h9225;
  rom[31069] = 16'h79e3;
  rom[31070] = 16'h9365;
  rom[31071] = 16'hf6cd;
  rom[31072] = 16'hff2a;
  rom[31073] = 16'hff0a;
  rom[31074] = 16'hff2b;
  rom[31075] = 16'hf72a;
  rom[31076] = 16'hff4a;
  rom[31077] = 16'hf749;
  rom[31078] = 16'hf74a;
  rom[31079] = 16'hef4a;
  rom[31080] = 16'hf74b;
  rom[31081] = 16'hf72a;
  rom[31082] = 16'hff49;
  rom[31083] = 16'hff28;
  rom[31084] = 16'hff48;
  rom[31085] = 16'hf748;
  rom[31086] = 16'hff69;
  rom[31087] = 16'hff4a;
  rom[31088] = 16'hf6ec;
  rom[31089] = 16'hf70d;
  rom[31090] = 16'hee6b;
  rom[31091] = 16'he5a9;
  rom[31092] = 16'hbc05;
  rom[31093] = 16'ha303;
  rom[31094] = 16'h8a01;
  rom[31095] = 16'h79a0;
  rom[31096] = 16'h81c1;
  rom[31097] = 16'h8a22;
  rom[31098] = 16'h81c1;
  rom[31099] = 16'h79e1;
  rom[31100] = 16'h8ac1;
  rom[31101] = 16'hbc45;
  rom[31102] = 16'hedc8;
  rom[31103] = 16'hfecc;
  rom[31104] = 16'hff2d;
  rom[31105] = 16'hf70b;
  rom[31106] = 16'he68a;
  rom[31107] = 16'ha4a5;
  rom[31108] = 16'h93e4;
  rom[31109] = 16'hcdca;
  rom[31110] = 16'hff4e;
  rom[31111] = 16'hf70a;
  rom[31112] = 16'hff4a;
  rom[31113] = 16'hf729;
  rom[31114] = 16'hff49;
  rom[31115] = 16'hf709;
  rom[31116] = 16'hff2a;
  rom[31117] = 16'hff09;
  rom[31118] = 16'hff2a;
  rom[31119] = 16'hff08;
  rom[31120] = 16'hff29;
  rom[31121] = 16'hff49;
  rom[31122] = 16'hff29;
  rom[31123] = 16'hff2a;
  rom[31124] = 16'hfeec;
  rom[31125] = 16'hbc86;
  rom[31126] = 16'ha263;
  rom[31127] = 16'hca66;
  rom[31128] = 16'hea47;
  rom[31129] = 16'hf226;
  rom[31130] = 16'hea67;
  rom[31131] = 16'hd267;
  rom[31132] = 16'hdb2b;
  rom[31133] = 16'hfd95;
  rom[31134] = 16'hff7d;
  rom[31135] = 16'hffde;
  rom[31136] = 16'hffff;
  rom[31137] = 16'hffff;
  rom[31138] = 16'hffff;
  rom[31139] = 16'hffff;
  rom[31140] = 16'hffff;
  rom[31141] = 16'hffff;
  rom[31142] = 16'hffff;
  rom[31143] = 16'hffff;
  rom[31144] = 16'hffff;
  rom[31145] = 16'hffff;
  rom[31146] = 16'hffff;
  rom[31147] = 16'hffff;
  rom[31148] = 16'hffff;
  rom[31149] = 16'hffff;
  rom[31150] = 16'hffff;
  rom[31151] = 16'hffff;
  rom[31152] = 16'hffff;
  rom[31153] = 16'hffff;
  rom[31154] = 16'hffff;
  rom[31155] = 16'hffff;
  rom[31156] = 16'hffff;
  rom[31157] = 16'hffff;
  rom[31158] = 16'hffff;
  rom[31159] = 16'hffff;
  rom[31160] = 16'hffff;
  rom[31161] = 16'hffff;
  rom[31162] = 16'hffff;
  rom[31163] = 16'hffff;
  rom[31164] = 16'hffff;
  rom[31165] = 16'hffff;
  rom[31166] = 16'hffff;
  rom[31167] = 16'hffff;
  rom[31168] = 16'hffff;
  rom[31169] = 16'hffff;
  rom[31170] = 16'hffff;
  rom[31171] = 16'hffff;
  rom[31172] = 16'hffff;
  rom[31173] = 16'hffff;
  rom[31174] = 16'hffff;
  rom[31175] = 16'hffff;
  rom[31176] = 16'hffff;
  rom[31177] = 16'hffff;
  rom[31178] = 16'hffff;
  rom[31179] = 16'hffff;
  rom[31180] = 16'hffff;
  rom[31181] = 16'hffff;
  rom[31182] = 16'hffff;
  rom[31183] = 16'hffff;
  rom[31184] = 16'hffff;
  rom[31185] = 16'hffff;
  rom[31186] = 16'hffff;
  rom[31187] = 16'hffff;
  rom[31188] = 16'hffff;
  rom[31189] = 16'hffff;
  rom[31190] = 16'hffff;
  rom[31191] = 16'hffff;
  rom[31192] = 16'hffff;
  rom[31193] = 16'hffff;
  rom[31194] = 16'hffff;
  rom[31195] = 16'hffff;
  rom[31196] = 16'hffff;
  rom[31197] = 16'hffff;
  rom[31198] = 16'hffff;
  rom[31199] = 16'hffff;
  rom[31200] = 16'hffff;
  rom[31201] = 16'hffff;
  rom[31202] = 16'hffff;
  rom[31203] = 16'hffff;
  rom[31204] = 16'hffff;
  rom[31205] = 16'hffff;
  rom[31206] = 16'hffff;
  rom[31207] = 16'hffff;
  rom[31208] = 16'hffff;
  rom[31209] = 16'hffff;
  rom[31210] = 16'hffff;
  rom[31211] = 16'hffff;
  rom[31212] = 16'hffff;
  rom[31213] = 16'hffff;
  rom[31214] = 16'hffff;
  rom[31215] = 16'hffdf;
  rom[31216] = 16'hffdf;
  rom[31217] = 16'hffde;
  rom[31218] = 16'hfeda;
  rom[31219] = 16'hf513;
  rom[31220] = 16'hca89;
  rom[31221] = 16'he249;
  rom[31222] = 16'hea07;
  rom[31223] = 16'hea47;
  rom[31224] = 16'he227;
  rom[31225] = 16'hea27;
  rom[31226] = 16'hea07;
  rom[31227] = 16'hf227;
  rom[31228] = 16'hea06;
  rom[31229] = 16'hf206;
  rom[31230] = 16'hf206;
  rom[31231] = 16'hea06;
  rom[31232] = 16'he206;
  rom[31233] = 16'hea26;
  rom[31234] = 16'hea06;
  rom[31235] = 16'hea27;
  rom[31236] = 16'he226;
  rom[31237] = 16'he206;
  rom[31238] = 16'hea06;
  rom[31239] = 16'hea28;
  rom[31240] = 16'hda48;
  rom[31241] = 16'ha9e4;
  rom[31242] = 16'ha2a3;
  rom[31243] = 16'he62c;
  rom[31244] = 16'heeeb;
  rom[31245] = 16'hf70b;
  rom[31246] = 16'hff0a;
  rom[31247] = 16'hff0a;
  rom[31248] = 16'hff29;
  rom[31249] = 16'hff29;
  rom[31250] = 16'hf708;
  rom[31251] = 16'hf74a;
  rom[31252] = 16'hef29;
  rom[31253] = 16'hf74a;
  rom[31254] = 16'hff0b;
  rom[31255] = 16'hff0c;
  rom[31256] = 16'hf6ca;
  rom[31257] = 16'hff2a;
  rom[31258] = 16'hf728;
  rom[31259] = 16'hf709;
  rom[31260] = 16'hf72a;
  rom[31261] = 16'hff0a;
  rom[31262] = 16'hef29;
  rom[31263] = 16'hef4a;
  rom[31264] = 16'hef2c;
  rom[31265] = 16'he60d;
  rom[31266] = 16'h8a83;
  rom[31267] = 16'ha204;
  rom[31268] = 16'hc266;
  rom[31269] = 16'h9a45;
  rom[31270] = 16'h8aa3;
  rom[31271] = 16'hf68c;
  rom[31272] = 16'hff09;
  rom[31273] = 16'hff29;
  rom[31274] = 16'hff09;
  rom[31275] = 16'hff29;
  rom[31276] = 16'hff07;
  rom[31277] = 16'hff28;
  rom[31278] = 16'hf728;
  rom[31279] = 16'hff2a;
  rom[31280] = 16'hf70a;
  rom[31281] = 16'hff2a;
  rom[31282] = 16'hf729;
  rom[31283] = 16'hff49;
  rom[31284] = 16'hf728;
  rom[31285] = 16'hff48;
  rom[31286] = 16'hf6c7;
  rom[31287] = 16'hff29;
  rom[31288] = 16'hf72a;
  rom[31289] = 16'hf72b;
  rom[31290] = 16'hf74b;
  rom[31291] = 16'hf6eb;
  rom[31292] = 16'hfecc;
  rom[31293] = 16'hee0a;
  rom[31294] = 16'hddea;
  rom[31295] = 16'hd5ca;
  rom[31296] = 16'hcd8a;
  rom[31297] = 16'hd56b;
  rom[31298] = 16'hdd8b;
  rom[31299] = 16'he60b;
  rom[31300] = 16'he689;
  rom[31301] = 16'hff2b;
  rom[31302] = 16'hf70a;
  rom[31303] = 16'hff2b;
  rom[31304] = 16'hf72c;
  rom[31305] = 16'he6cc;
  rom[31306] = 16'h9ca5;
  rom[31307] = 16'h8c03;
  rom[31308] = 16'hde6b;
  rom[31309] = 16'hf70c;
  rom[31310] = 16'hf709;
  rom[31311] = 16'hf749;
  rom[31312] = 16'hef27;
  rom[31313] = 16'hf72a;
  rom[31314] = 16'hf709;
  rom[31315] = 16'hff0a;
  rom[31316] = 16'hf70a;
  rom[31317] = 16'hff0a;
  rom[31318] = 16'hff0a;
  rom[31319] = 16'hff0a;
  rom[31320] = 16'hf70a;
  rom[31321] = 16'hff29;
  rom[31322] = 16'hf6e8;
  rom[31323] = 16'hff4a;
  rom[31324] = 16'hf70b;
  rom[31325] = 16'hcd69;
  rom[31326] = 16'h92a4;
  rom[31327] = 16'hca88;
  rom[31328] = 16'he206;
  rom[31329] = 16'hf207;
  rom[31330] = 16'he227;
  rom[31331] = 16'hca89;
  rom[31332] = 16'hdc70;
  rom[31333] = 16'hff1a;
  rom[31334] = 16'hffbe;
  rom[31335] = 16'hffff;
  rom[31336] = 16'hffff;
  rom[31337] = 16'hffff;
  rom[31338] = 16'hffff;
  rom[31339] = 16'hffff;
  rom[31340] = 16'hffff;
  rom[31341] = 16'hf7ff;
  rom[31342] = 16'hf7ff;
  rom[31343] = 16'hffff;
  rom[31344] = 16'hffff;
  rom[31345] = 16'hffff;
  rom[31346] = 16'hffff;
  rom[31347] = 16'hffff;
  rom[31348] = 16'hffff;
  rom[31349] = 16'hffff;
  rom[31350] = 16'hffff;
  rom[31351] = 16'hffff;
  rom[31352] = 16'hffff;
  rom[31353] = 16'hffff;
  rom[31354] = 16'hffff;
  rom[31355] = 16'hffff;
  rom[31356] = 16'hffff;
  rom[31357] = 16'hffff;
  rom[31358] = 16'hffff;
  rom[31359] = 16'hffff;
  rom[31360] = 16'hffff;
  rom[31361] = 16'hffff;
  rom[31362] = 16'hfffe;
  rom[31363] = 16'hffff;
  rom[31364] = 16'hffff;
  rom[31365] = 16'hffff;
  rom[31366] = 16'hffff;
  rom[31367] = 16'hffff;
  rom[31368] = 16'hffff;
  rom[31369] = 16'hffff;
  rom[31370] = 16'hffff;
  rom[31371] = 16'hffff;
  rom[31372] = 16'hffff;
  rom[31373] = 16'hffff;
  rom[31374] = 16'hffff;
  rom[31375] = 16'hffff;
  rom[31376] = 16'hffff;
  rom[31377] = 16'hffff;
  rom[31378] = 16'hffff;
  rom[31379] = 16'hffff;
  rom[31380] = 16'hffff;
  rom[31381] = 16'hffff;
  rom[31382] = 16'hffff;
  rom[31383] = 16'hffff;
  rom[31384] = 16'hffff;
  rom[31385] = 16'hffff;
  rom[31386] = 16'hffff;
  rom[31387] = 16'hffff;
  rom[31388] = 16'hffff;
  rom[31389] = 16'hffff;
  rom[31390] = 16'hffff;
  rom[31391] = 16'hffff;
  rom[31392] = 16'hffff;
  rom[31393] = 16'hffff;
  rom[31394] = 16'hffff;
  rom[31395] = 16'hffff;
  rom[31396] = 16'hffff;
  rom[31397] = 16'hffff;
  rom[31398] = 16'hffff;
  rom[31399] = 16'hffff;
  rom[31400] = 16'hffff;
  rom[31401] = 16'hffff;
  rom[31402] = 16'hffff;
  rom[31403] = 16'hffff;
  rom[31404] = 16'hffff;
  rom[31405] = 16'hffff;
  rom[31406] = 16'hffff;
  rom[31407] = 16'hffff;
  rom[31408] = 16'hffff;
  rom[31409] = 16'hffff;
  rom[31410] = 16'hffff;
  rom[31411] = 16'hffff;
  rom[31412] = 16'hffff;
  rom[31413] = 16'hffff;
  rom[31414] = 16'hffff;
  rom[31415] = 16'hffff;
  rom[31416] = 16'hffff;
  rom[31417] = 16'hffff;
  rom[31418] = 16'hffde;
  rom[31419] = 16'hff1b;
  rom[31420] = 16'hf4f3;
  rom[31421] = 16'hc269;
  rom[31422] = 16'he28a;
  rom[31423] = 16'hda27;
  rom[31424] = 16'he267;
  rom[31425] = 16'hea27;
  rom[31426] = 16'hf248;
  rom[31427] = 16'hea06;
  rom[31428] = 16'hf226;
  rom[31429] = 16'hf206;
  rom[31430] = 16'hf227;
  rom[31431] = 16'hf207;
  rom[31432] = 16'hea46;
  rom[31433] = 16'hea26;
  rom[31434] = 16'hf227;
  rom[31435] = 16'hea06;
  rom[31436] = 16'hea47;
  rom[31437] = 16'he226;
  rom[31438] = 16'hea28;
  rom[31439] = 16'hea27;
  rom[31440] = 16'hea49;
  rom[31441] = 16'hd247;
  rom[31442] = 16'h9182;
  rom[31443] = 16'h9302;
  rom[31444] = 16'hee8d;
  rom[31445] = 16'hff0c;
  rom[31446] = 16'hf6aa;
  rom[31447] = 16'hfeea;
  rom[31448] = 16'hff0a;
  rom[31449] = 16'hff29;
  rom[31450] = 16'hff2a;
  rom[31451] = 16'hf749;
  rom[31452] = 16'hf769;
  rom[31453] = 16'hef07;
  rom[31454] = 16'hff09;
  rom[31455] = 16'hff2a;
  rom[31456] = 16'hff2a;
  rom[31457] = 16'hf729;
  rom[31458] = 16'hff8a;
  rom[31459] = 16'hff49;
  rom[31460] = 16'hff4a;
  rom[31461] = 16'hf74a;
  rom[31462] = 16'hef2b;
  rom[31463] = 16'hf74c;
  rom[31464] = 16'hf6ae;
  rom[31465] = 16'h8a41;
  rom[31466] = 16'h99e4;
  rom[31467] = 16'hd267;
  rom[31468] = 16'he287;
  rom[31469] = 16'haa05;
  rom[31470] = 16'h8a42;
  rom[31471] = 16'hedea;
  rom[31472] = 16'hff4a;
  rom[31473] = 16'hf708;
  rom[31474] = 16'hff2a;
  rom[31475] = 16'hff29;
  rom[31476] = 16'hff28;
  rom[31477] = 16'hff27;
  rom[31478] = 16'hff08;
  rom[31479] = 16'hff09;
  rom[31480] = 16'hff2a;
  rom[31481] = 16'hff29;
  rom[31482] = 16'hff2a;
  rom[31483] = 16'hff09;
  rom[31484] = 16'hff29;
  rom[31485] = 16'hff28;
  rom[31486] = 16'hff4a;
  rom[31487] = 16'hff29;
  rom[31488] = 16'heee8;
  rom[31489] = 16'hf748;
  rom[31490] = 16'hff6a;
  rom[31491] = 16'hff4a;
  rom[31492] = 16'hff0b;
  rom[31493] = 16'hfeea;
  rom[31494] = 16'heeea;
  rom[31495] = 16'hf72b;
  rom[31496] = 16'hf72c;
  rom[31497] = 16'hf72d;
  rom[31498] = 16'hff0d;
  rom[31499] = 16'hf6eb;
  rom[31500] = 16'heee9;
  rom[31501] = 16'hf729;
  rom[31502] = 16'hff8b;
  rom[31503] = 16'hef0a;
  rom[31504] = 16'hffaf;
  rom[31505] = 16'h9c65;
  rom[31506] = 16'h83a5;
  rom[31507] = 16'he6cd;
  rom[31508] = 16'hff2c;
  rom[31509] = 16'hf708;
  rom[31510] = 16'hff49;
  rom[31511] = 16'hff67;
  rom[31512] = 16'hf747;
  rom[31513] = 16'hf729;
  rom[31514] = 16'hf70a;
  rom[31515] = 16'hff2a;
  rom[31516] = 16'hf6ea;
  rom[31517] = 16'hff0a;
  rom[31518] = 16'hff2a;
  rom[31519] = 16'hff2a;
  rom[31520] = 16'hff2a;
  rom[31521] = 16'hff4a;
  rom[31522] = 16'hff2a;
  rom[31523] = 16'hf709;
  rom[31524] = 16'hf72b;
  rom[31525] = 16'hde0c;
  rom[31526] = 16'hab88;
  rom[31527] = 16'hca88;
  rom[31528] = 16'hea08;
  rom[31529] = 16'hf207;
  rom[31530] = 16'he248;
  rom[31531] = 16'hc2c9;
  rom[31532] = 16'hfe58;
  rom[31533] = 16'hff9c;
  rom[31534] = 16'hffff;
  rom[31535] = 16'hffff;
  rom[31536] = 16'hffff;
  rom[31537] = 16'hffff;
  rom[31538] = 16'hffff;
  rom[31539] = 16'hffff;
  rom[31540] = 16'hffff;
  rom[31541] = 16'hffff;
  rom[31542] = 16'hffff;
  rom[31543] = 16'hffff;
  rom[31544] = 16'hffff;
  rom[31545] = 16'hffff;
  rom[31546] = 16'hffff;
  rom[31547] = 16'hffff;
  rom[31548] = 16'hffff;
  rom[31549] = 16'hffff;
  rom[31550] = 16'hffff;
  rom[31551] = 16'hffff;
  rom[31552] = 16'hffff;
  rom[31553] = 16'hffff;
  rom[31554] = 16'hffff;
  rom[31555] = 16'hffff;
  rom[31556] = 16'hffff;
  rom[31557] = 16'hffff;
  rom[31558] = 16'hffff;
  rom[31559] = 16'hffff;
  rom[31560] = 16'hffff;
  rom[31561] = 16'hffff;
  rom[31562] = 16'hffff;
  rom[31563] = 16'hffff;
  rom[31564] = 16'hffff;
  rom[31565] = 16'hffff;
  rom[31566] = 16'hffff;
  rom[31567] = 16'hffff;
  rom[31568] = 16'hffff;
  rom[31569] = 16'hffff;
  rom[31570] = 16'hffff;
  rom[31571] = 16'hffff;
  rom[31572] = 16'hffff;
  rom[31573] = 16'hffff;
  rom[31574] = 16'hffff;
  rom[31575] = 16'hffff;
  rom[31576] = 16'hffff;
  rom[31577] = 16'hffff;
  rom[31578] = 16'hffff;
  rom[31579] = 16'hffff;
  rom[31580] = 16'hffff;
  rom[31581] = 16'hffff;
  rom[31582] = 16'hffff;
  rom[31583] = 16'hffff;
  rom[31584] = 16'hffff;
  rom[31585] = 16'hffff;
  rom[31586] = 16'hffff;
  rom[31587] = 16'hffff;
  rom[31588] = 16'hffff;
  rom[31589] = 16'hffff;
  rom[31590] = 16'hffff;
  rom[31591] = 16'hffff;
  rom[31592] = 16'hffff;
  rom[31593] = 16'hffff;
  rom[31594] = 16'hffff;
  rom[31595] = 16'hffff;
  rom[31596] = 16'hffff;
  rom[31597] = 16'hffff;
  rom[31598] = 16'hffff;
  rom[31599] = 16'hffff;
  rom[31600] = 16'hffff;
  rom[31601] = 16'hffff;
  rom[31602] = 16'hffff;
  rom[31603] = 16'hffff;
  rom[31604] = 16'hffff;
  rom[31605] = 16'hffff;
  rom[31606] = 16'hffff;
  rom[31607] = 16'hffff;
  rom[31608] = 16'hffff;
  rom[31609] = 16'hffff;
  rom[31610] = 16'hffff;
  rom[31611] = 16'hffff;
  rom[31612] = 16'hffff;
  rom[31613] = 16'hffff;
  rom[31614] = 16'hfffe;
  rom[31615] = 16'hffff;
  rom[31616] = 16'hffff;
  rom[31617] = 16'hffff;
  rom[31618] = 16'hffff;
  rom[31619] = 16'hffbe;
  rom[31620] = 16'hfefa;
  rom[31621] = 16'hed54;
  rom[31622] = 16'hc32b;
  rom[31623] = 16'hd289;
  rom[31624] = 16'hda27;
  rom[31625] = 16'hea28;
  rom[31626] = 16'hea27;
  rom[31627] = 16'he227;
  rom[31628] = 16'hea26;
  rom[31629] = 16'hf207;
  rom[31630] = 16'hf207;
  rom[31631] = 16'hf207;
  rom[31632] = 16'hea07;
  rom[31633] = 16'hea47;
  rom[31634] = 16'hea06;
  rom[31635] = 16'hea06;
  rom[31636] = 16'hea26;
  rom[31637] = 16'hea47;
  rom[31638] = 16'he207;
  rom[31639] = 16'hf1e7;
  rom[31640] = 16'he9e7;
  rom[31641] = 16'he226;
  rom[31642] = 16'hc265;
  rom[31643] = 16'h81e1;
  rom[31644] = 16'h9344;
  rom[31645] = 16'hee0b;
  rom[31646] = 16'hfeec;
  rom[31647] = 16'hfeeb;
  rom[31648] = 16'hf6ea;
  rom[31649] = 16'hff4a;
  rom[31650] = 16'hf708;
  rom[31651] = 16'hff28;
  rom[31652] = 16'hff08;
  rom[31653] = 16'hff08;
  rom[31654] = 16'hff08;
  rom[31655] = 16'hff09;
  rom[31656] = 16'hf709;
  rom[31657] = 16'hff4b;
  rom[31658] = 16'hf6e9;
  rom[31659] = 16'hff2b;
  rom[31660] = 16'hf70a;
  rom[31661] = 16'hf72b;
  rom[31662] = 16'hf74d;
  rom[31663] = 16'he60b;
  rom[31664] = 16'h8a61;
  rom[31665] = 16'h99c3;
  rom[31666] = 16'hca67;
  rom[31667] = 16'hda48;
  rom[31668] = 16'hda46;
  rom[31669] = 16'hba66;
  rom[31670] = 16'h89e1;
  rom[31671] = 16'hdd49;
  rom[31672] = 16'hff0a;
  rom[31673] = 16'hf729;
  rom[31674] = 16'hf729;
  rom[31675] = 16'hf72a;
  rom[31676] = 16'hf708;
  rom[31677] = 16'hff29;
  rom[31678] = 16'hff08;
  rom[31679] = 16'hff08;
  rom[31680] = 16'hff09;
  rom[31681] = 16'hff09;
  rom[31682] = 16'hf709;
  rom[31683] = 16'hff29;
  rom[31684] = 16'hff09;
  rom[31685] = 16'hff29;
  rom[31686] = 16'hf708;
  rom[31687] = 16'hf709;
  rom[31688] = 16'hf708;
  rom[31689] = 16'hf74a;
  rom[31690] = 16'hf729;
  rom[31691] = 16'hff0a;
  rom[31692] = 16'hff09;
  rom[31693] = 16'hff2a;
  rom[31694] = 16'hff0a;
  rom[31695] = 16'hff0a;
  rom[31696] = 16'hff09;
  rom[31697] = 16'hff0a;
  rom[31698] = 16'hf709;
  rom[31699] = 16'hff4b;
  rom[31700] = 16'hf728;
  rom[31701] = 16'hf729;
  rom[31702] = 16'hef0a;
  rom[31703] = 16'hf72d;
  rom[31704] = 16'hb4e7;
  rom[31705] = 16'h7b42;
  rom[31706] = 16'hce0a;
  rom[31707] = 16'hf72d;
  rom[31708] = 16'heee9;
  rom[31709] = 16'hf729;
  rom[31710] = 16'hf728;
  rom[31711] = 16'hf728;
  rom[31712] = 16'hff28;
  rom[31713] = 16'hff29;
  rom[31714] = 16'hf708;
  rom[31715] = 16'hff08;
  rom[31716] = 16'hff08;
  rom[31717] = 16'hff29;
  rom[31718] = 16'hef28;
  rom[31719] = 16'hf729;
  rom[31720] = 16'hf708;
  rom[31721] = 16'hff29;
  rom[31722] = 16'hf709;
  rom[31723] = 16'hf72a;
  rom[31724] = 16'hf6ea;
  rom[31725] = 16'he64d;
  rom[31726] = 16'hab88;
  rom[31727] = 16'hcaa8;
  rom[31728] = 16'he9e6;
  rom[31729] = 16'hf9e8;
  rom[31730] = 16'hd249;
  rom[31731] = 16'hcbce;
  rom[31732] = 16'hff5b;
  rom[31733] = 16'hffdd;
  rom[31734] = 16'hffff;
  rom[31735] = 16'hffff;
  rom[31736] = 16'hffff;
  rom[31737] = 16'hffff;
  rom[31738] = 16'hffff;
  rom[31739] = 16'hffff;
  rom[31740] = 16'hffff;
  rom[31741] = 16'hffff;
  rom[31742] = 16'hffff;
  rom[31743] = 16'hffff;
  rom[31744] = 16'hffff;
  rom[31745] = 16'hffff;
  rom[31746] = 16'hffff;
  rom[31747] = 16'hffff;
  rom[31748] = 16'hffff;
  rom[31749] = 16'hffff;
  rom[31750] = 16'hffff;
  rom[31751] = 16'hffff;
  rom[31752] = 16'hffff;
  rom[31753] = 16'hffff;
  rom[31754] = 16'hffff;
  rom[31755] = 16'hffff;
  rom[31756] = 16'hffff;
  rom[31757] = 16'hffff;
  rom[31758] = 16'hffff;
  rom[31759] = 16'hffff;
  rom[31760] = 16'hffff;
  rom[31761] = 16'hffff;
  rom[31762] = 16'hffff;
  rom[31763] = 16'hffff;
  rom[31764] = 16'hffff;
  rom[31765] = 16'hffff;
  rom[31766] = 16'hffff;
  rom[31767] = 16'hffff;
  rom[31768] = 16'hffff;
  rom[31769] = 16'hffff;
  rom[31770] = 16'hffff;
  rom[31771] = 16'hffff;
  rom[31772] = 16'hffff;
  rom[31773] = 16'hffff;
  rom[31774] = 16'hffff;
  rom[31775] = 16'hffff;
  rom[31776] = 16'hffff;
  rom[31777] = 16'hffff;
  rom[31778] = 16'hffff;
  rom[31779] = 16'hffff;
  rom[31780] = 16'hffff;
  rom[31781] = 16'hffff;
  rom[31782] = 16'hffff;
  rom[31783] = 16'hffff;
  rom[31784] = 16'hffff;
  rom[31785] = 16'hffff;
  rom[31786] = 16'hffff;
  rom[31787] = 16'hffff;
  rom[31788] = 16'hffff;
  rom[31789] = 16'hffff;
  rom[31790] = 16'hffff;
  rom[31791] = 16'hffff;
  rom[31792] = 16'hffff;
  rom[31793] = 16'hffff;
  rom[31794] = 16'hffff;
  rom[31795] = 16'hffff;
  rom[31796] = 16'hffff;
  rom[31797] = 16'hffff;
  rom[31798] = 16'hffff;
  rom[31799] = 16'hffff;
  rom[31800] = 16'hffff;
  rom[31801] = 16'hffff;
  rom[31802] = 16'hffff;
  rom[31803] = 16'hffff;
  rom[31804] = 16'hffff;
  rom[31805] = 16'hffff;
  rom[31806] = 16'hffff;
  rom[31807] = 16'hffff;
  rom[31808] = 16'hffff;
  rom[31809] = 16'hffff;
  rom[31810] = 16'hffff;
  rom[31811] = 16'hffff;
  rom[31812] = 16'hffff;
  rom[31813] = 16'hffff;
  rom[31814] = 16'hffff;
  rom[31815] = 16'hffff;
  rom[31816] = 16'hffff;
  rom[31817] = 16'hffff;
  rom[31818] = 16'hffff;
  rom[31819] = 16'hffdf;
  rom[31820] = 16'hffdf;
  rom[31821] = 16'hff3b;
  rom[31822] = 16'hfdd7;
  rom[31823] = 16'hd38d;
  rom[31824] = 16'hd289;
  rom[31825] = 16'he268;
  rom[31826] = 16'he247;
  rom[31827] = 16'he246;
  rom[31828] = 16'hea26;
  rom[31829] = 16'hf226;
  rom[31830] = 16'hf1e6;
  rom[31831] = 16'hf1e6;
  rom[31832] = 16'hf207;
  rom[31833] = 16'hf206;
  rom[31834] = 16'hf226;
  rom[31835] = 16'hea26;
  rom[31836] = 16'hea27;
  rom[31837] = 16'he206;
  rom[31838] = 16'hea27;
  rom[31839] = 16'hea07;
  rom[31840] = 16'hf207;
  rom[31841] = 16'hea47;
  rom[31842] = 16'hd247;
  rom[31843] = 16'hbac6;
  rom[31844] = 16'h8a23;
  rom[31845] = 16'h8ac2;
  rom[31846] = 16'he58b;
  rom[31847] = 16'hfeee;
  rom[31848] = 16'hf70c;
  rom[31849] = 16'hf72b;
  rom[31850] = 16'hf729;
  rom[31851] = 16'hf728;
  rom[31852] = 16'hff07;
  rom[31853] = 16'hff28;
  rom[31854] = 16'hff08;
  rom[31855] = 16'hff08;
  rom[31856] = 16'hff29;
  rom[31857] = 16'hff29;
  rom[31858] = 16'hff0a;
  rom[31859] = 16'hfeea;
  rom[31860] = 16'hff2d;
  rom[31861] = 16'hf70e;
  rom[31862] = 16'hddcb;
  rom[31863] = 16'h92a3;
  rom[31864] = 16'hb265;
  rom[31865] = 16'hca06;
  rom[31866] = 16'hea69;
  rom[31867] = 16'he1e7;
  rom[31868] = 16'he268;
  rom[31869] = 16'hcaa8;
  rom[31870] = 16'h89c2;
  rom[31871] = 16'hbc67;
  rom[31872] = 16'hff2b;
  rom[31873] = 16'hf709;
  rom[31874] = 16'hff6a;
  rom[31875] = 16'hf72a;
  rom[31876] = 16'hf72a;
  rom[31877] = 16'hff29;
  rom[31878] = 16'hff29;
  rom[31879] = 16'hff28;
  rom[31880] = 16'hff29;
  rom[31881] = 16'hff09;
  rom[31882] = 16'hff2a;
  rom[31883] = 16'hff29;
  rom[31884] = 16'hff2a;
  rom[31885] = 16'hff09;
  rom[31886] = 16'hf709;
  rom[31887] = 16'hf729;
  rom[31888] = 16'hff4a;
  rom[31889] = 16'hf728;
  rom[31890] = 16'hff2a;
  rom[31891] = 16'hfee9;
  rom[31892] = 16'hff29;
  rom[31893] = 16'hff29;
  rom[31894] = 16'hff2a;
  rom[31895] = 16'hff09;
  rom[31896] = 16'hff29;
  rom[31897] = 16'hff09;
  rom[31898] = 16'hff2a;
  rom[31899] = 16'hf709;
  rom[31900] = 16'hff69;
  rom[31901] = 16'hf74a;
  rom[31902] = 16'hf72d;
  rom[31903] = 16'hd62b;
  rom[31904] = 16'h7b41;
  rom[31905] = 16'hd5ea;
  rom[31906] = 16'hff2d;
  rom[31907] = 16'hf72a;
  rom[31908] = 16'hff6a;
  rom[31909] = 16'hff6a;
  rom[31910] = 16'hff6a;
  rom[31911] = 16'hf708;
  rom[31912] = 16'hff49;
  rom[31913] = 16'hff28;
  rom[31914] = 16'hff09;
  rom[31915] = 16'hff08;
  rom[31916] = 16'hff29;
  rom[31917] = 16'hf728;
  rom[31918] = 16'hf749;
  rom[31919] = 16'hf729;
  rom[31920] = 16'hff4a;
  rom[31921] = 16'hfee9;
  rom[31922] = 16'hff2a;
  rom[31923] = 16'hf72a;
  rom[31924] = 16'hff2c;
  rom[31925] = 16'hddec;
  rom[31926] = 16'ha367;
  rom[31927] = 16'hc287;
  rom[31928] = 16'hf207;
  rom[31929] = 16'hf207;
  rom[31930] = 16'hca69;
  rom[31931] = 16'hed54;
  rom[31932] = 16'hffbd;
  rom[31933] = 16'hfffe;
  rom[31934] = 16'hffff;
  rom[31935] = 16'hffdf;
  rom[31936] = 16'hffdf;
  rom[31937] = 16'hffff;
  rom[31938] = 16'hffff;
  rom[31939] = 16'hffff;
  rom[31940] = 16'hffff;
  rom[31941] = 16'hffff;
  rom[31942] = 16'hffff;
  rom[31943] = 16'hffff;
  rom[31944] = 16'hffff;
  rom[31945] = 16'hffff;
  rom[31946] = 16'hffff;
  rom[31947] = 16'hffff;
  rom[31948] = 16'hffff;
  rom[31949] = 16'hffff;
  rom[31950] = 16'hffff;
  rom[31951] = 16'hffff;
  rom[31952] = 16'hffff;
  rom[31953] = 16'hffff;
  rom[31954] = 16'hffff;
  rom[31955] = 16'hffff;
  rom[31956] = 16'hffff;
  rom[31957] = 16'hffff;
  rom[31958] = 16'hffff;
  rom[31959] = 16'hffff;
  rom[31960] = 16'hffff;
  rom[31961] = 16'hffff;
  rom[31962] = 16'hffff;
  rom[31963] = 16'hffff;
  rom[31964] = 16'hffff;
  rom[31965] = 16'hffff;
  rom[31966] = 16'hffff;
  rom[31967] = 16'hffff;
  rom[31968] = 16'hffff;
  rom[31969] = 16'hffff;
  rom[31970] = 16'hffff;
  rom[31971] = 16'hffff;
  rom[31972] = 16'hffff;
  rom[31973] = 16'hffff;
  rom[31974] = 16'hffff;
  rom[31975] = 16'hffff;
  rom[31976] = 16'hffff;
  rom[31977] = 16'hffff;
  rom[31978] = 16'hffff;
  rom[31979] = 16'hffff;
  rom[31980] = 16'hffff;
  rom[31981] = 16'hffff;
  rom[31982] = 16'hffff;
  rom[31983] = 16'hffff;
  rom[31984] = 16'hffff;
  rom[31985] = 16'hffff;
  rom[31986] = 16'hffff;
  rom[31987] = 16'hffff;
  rom[31988] = 16'hffff;
  rom[31989] = 16'hffff;
  rom[31990] = 16'hffff;
  rom[31991] = 16'hffff;
  rom[31992] = 16'hffff;
  rom[31993] = 16'hffff;
  rom[31994] = 16'hffff;
  rom[31995] = 16'hffff;
  rom[31996] = 16'hffff;
  rom[31997] = 16'hffff;
  rom[31998] = 16'hffff;
  rom[31999] = 16'hffff;
  rom[32000] = 16'hffff;
  rom[32001] = 16'hffff;
  rom[32002] = 16'hffff;
  rom[32003] = 16'hffff;
  rom[32004] = 16'hffff;
  rom[32005] = 16'hffff;
  rom[32006] = 16'hffff;
  rom[32007] = 16'hffff;
  rom[32008] = 16'hffff;
  rom[32009] = 16'hffff;
  rom[32010] = 16'hffff;
  rom[32011] = 16'hffff;
  rom[32012] = 16'hffff;
  rom[32013] = 16'hffff;
  rom[32014] = 16'hffff;
  rom[32015] = 16'hffff;
  rom[32016] = 16'hffff;
  rom[32017] = 16'hffff;
  rom[32018] = 16'hffff;
  rom[32019] = 16'hffff;
  rom[32020] = 16'hffdf;
  rom[32021] = 16'hfffe;
  rom[32022] = 16'hff7d;
  rom[32023] = 16'hfeda;
  rom[32024] = 16'hecd1;
  rom[32025] = 16'hcb0a;
  rom[32026] = 16'hd2c8;
  rom[32027] = 16'hd266;
  rom[32028] = 16'hda45;
  rom[32029] = 16'hea46;
  rom[32030] = 16'hf206;
  rom[32031] = 16'hfa06;
  rom[32032] = 16'hf206;
  rom[32033] = 16'hf1e6;
  rom[32034] = 16'hf206;
  rom[32035] = 16'hf226;
  rom[32036] = 16'he226;
  rom[32037] = 16'hea47;
  rom[32038] = 16'hea27;
  rom[32039] = 16'hf227;
  rom[32040] = 16'hf227;
  rom[32041] = 16'hea07;
  rom[32042] = 16'he247;
  rom[32043] = 16'hca87;
  rom[32044] = 16'hb286;
  rom[32045] = 16'h9223;
  rom[32046] = 16'h7a02;
  rom[32047] = 16'hbc48;
  rom[32048] = 16'hf68d;
  rom[32049] = 16'hf6ed;
  rom[32050] = 16'hf72b;
  rom[32051] = 16'hf72a;
  rom[32052] = 16'hf728;
  rom[32053] = 16'hff49;
  rom[32054] = 16'hff29;
  rom[32055] = 16'hff49;
  rom[32056] = 16'hf709;
  rom[32057] = 16'hff4a;
  rom[32058] = 16'hfeeb;
  rom[32059] = 16'hff0d;
  rom[32060] = 16'hf68d;
  rom[32061] = 16'hd52b;
  rom[32062] = 16'h9283;
  rom[32063] = 16'h99c4;
  rom[32064] = 16'hca05;
  rom[32065] = 16'hea28;
  rom[32066] = 16'hf1e7;
  rom[32067] = 16'hfa48;
  rom[32068] = 16'he206;
  rom[32069] = 16'hd268;
  rom[32070] = 16'h89c3;
  rom[32071] = 16'h9b64;
  rom[32072] = 16'hff0d;
  rom[32073] = 16'hf6c9;
  rom[32074] = 16'hff6a;
  rom[32075] = 16'hf749;
  rom[32076] = 16'hef09;
  rom[32077] = 16'hf749;
  rom[32078] = 16'hf709;
  rom[32079] = 16'hff28;
  rom[32080] = 16'hf708;
  rom[32081] = 16'hff29;
  rom[32082] = 16'hff09;
  rom[32083] = 16'hff29;
  rom[32084] = 16'hf709;
  rom[32085] = 16'hff29;
  rom[32086] = 16'hff29;
  rom[32087] = 16'hff29;
  rom[32088] = 16'hef09;
  rom[32089] = 16'hf729;
  rom[32090] = 16'hff09;
  rom[32091] = 16'hff29;
  rom[32092] = 16'hf708;
  rom[32093] = 16'hff29;
  rom[32094] = 16'hff29;
  rom[32095] = 16'hff09;
  rom[32096] = 16'hf6e8;
  rom[32097] = 16'hf6e8;
  rom[32098] = 16'hff29;
  rom[32099] = 16'hf749;
  rom[32100] = 16'hef08;
  rom[32101] = 16'hf72b;
  rom[32102] = 16'heeee;
  rom[32103] = 16'h8ba3;
  rom[32104] = 16'hb508;
  rom[32105] = 16'heecc;
  rom[32106] = 16'hff4b;
  rom[32107] = 16'heee8;
  rom[32108] = 16'hf768;
  rom[32109] = 16'hf728;
  rom[32110] = 16'hf709;
  rom[32111] = 16'hff09;
  rom[32112] = 16'hf708;
  rom[32113] = 16'hff28;
  rom[32114] = 16'hfee9;
  rom[32115] = 16'hff09;
  rom[32116] = 16'hf709;
  rom[32117] = 16'hf749;
  rom[32118] = 16'hf729;
  rom[32119] = 16'hff29;
  rom[32120] = 16'hff0a;
  rom[32121] = 16'hfeca;
  rom[32122] = 16'hff0a;
  rom[32123] = 16'hff0b;
  rom[32124] = 16'hfeea;
  rom[32125] = 16'hddcb;
  rom[32126] = 16'h92a4;
  rom[32127] = 16'hcaa7;
  rom[32128] = 16'hea26;
  rom[32129] = 16'hea47;
  rom[32130] = 16'hcaca;
  rom[32131] = 16'hfedb;
  rom[32132] = 16'hffbd;
  rom[32133] = 16'hffff;
  rom[32134] = 16'hffff;
  rom[32135] = 16'hffff;
  rom[32136] = 16'hffff;
  rom[32137] = 16'hffff;
  rom[32138] = 16'hffff;
  rom[32139] = 16'hffff;
  rom[32140] = 16'hffff;
  rom[32141] = 16'hffff;
  rom[32142] = 16'hffff;
  rom[32143] = 16'hffff;
  rom[32144] = 16'hffff;
  rom[32145] = 16'hffff;
  rom[32146] = 16'hffff;
  rom[32147] = 16'hffff;
  rom[32148] = 16'hffff;
  rom[32149] = 16'hffff;
  rom[32150] = 16'hffff;
  rom[32151] = 16'hffff;
  rom[32152] = 16'hffff;
  rom[32153] = 16'hffff;
  rom[32154] = 16'hffff;
  rom[32155] = 16'hffff;
  rom[32156] = 16'hffff;
  rom[32157] = 16'hffff;
  rom[32158] = 16'hffff;
  rom[32159] = 16'hffff;
  rom[32160] = 16'hffff;
  rom[32161] = 16'hffff;
  rom[32162] = 16'hffff;
  rom[32163] = 16'hffff;
  rom[32164] = 16'hffff;
  rom[32165] = 16'hffff;
  rom[32166] = 16'hffff;
  rom[32167] = 16'hffff;
  rom[32168] = 16'hffff;
  rom[32169] = 16'hffff;
  rom[32170] = 16'hffff;
  rom[32171] = 16'hffff;
  rom[32172] = 16'hffff;
  rom[32173] = 16'hffff;
  rom[32174] = 16'hffff;
  rom[32175] = 16'hffff;
  rom[32176] = 16'hffff;
  rom[32177] = 16'hffff;
  rom[32178] = 16'hffff;
  rom[32179] = 16'hffff;
  rom[32180] = 16'hffff;
  rom[32181] = 16'hffff;
  rom[32182] = 16'hffff;
  rom[32183] = 16'hffff;
  rom[32184] = 16'hffff;
  rom[32185] = 16'hffff;
  rom[32186] = 16'hffff;
  rom[32187] = 16'hffff;
  rom[32188] = 16'hffff;
  rom[32189] = 16'hffff;
  rom[32190] = 16'hffff;
  rom[32191] = 16'hffff;
  rom[32192] = 16'hffff;
  rom[32193] = 16'hffff;
  rom[32194] = 16'hffff;
  rom[32195] = 16'hffff;
  rom[32196] = 16'hffff;
  rom[32197] = 16'hffff;
  rom[32198] = 16'hffff;
  rom[32199] = 16'hffff;
  rom[32200] = 16'hffff;
  rom[32201] = 16'hffff;
  rom[32202] = 16'hffff;
  rom[32203] = 16'hffff;
  rom[32204] = 16'hffff;
  rom[32205] = 16'hffff;
  rom[32206] = 16'hffff;
  rom[32207] = 16'hffff;
  rom[32208] = 16'hffff;
  rom[32209] = 16'hffff;
  rom[32210] = 16'hffff;
  rom[32211] = 16'hffff;
  rom[32212] = 16'hffff;
  rom[32213] = 16'hffff;
  rom[32214] = 16'hffff;
  rom[32215] = 16'hffff;
  rom[32216] = 16'hffff;
  rom[32217] = 16'hffff;
  rom[32218] = 16'hffff;
  rom[32219] = 16'hffff;
  rom[32220] = 16'hffff;
  rom[32221] = 16'hffff;
  rom[32222] = 16'hffff;
  rom[32223] = 16'hffbd;
  rom[32224] = 16'hff5c;
  rom[32225] = 16'hfe57;
  rom[32226] = 16'hed12;
  rom[32227] = 16'hcb2a;
  rom[32228] = 16'hc267;
  rom[32229] = 16'hdaa8;
  rom[32230] = 16'he228;
  rom[32231] = 16'hea07;
  rom[32232] = 16'hf227;
  rom[32233] = 16'hea06;
  rom[32234] = 16'hf227;
  rom[32235] = 16'hea26;
  rom[32236] = 16'hf267;
  rom[32237] = 16'hea47;
  rom[32238] = 16'hea47;
  rom[32239] = 16'hea07;
  rom[32240] = 16'hf207;
  rom[32241] = 16'hea07;
  rom[32242] = 16'hea28;
  rom[32243] = 16'he248;
  rom[32244] = 16'hda88;
  rom[32245] = 16'hc266;
  rom[32246] = 16'haa65;
  rom[32247] = 16'h89e2;
  rom[32248] = 16'h8a63;
  rom[32249] = 16'hbc67;
  rom[32250] = 16'hf6cf;
  rom[32251] = 16'hff0e;
  rom[32252] = 16'hff0d;
  rom[32253] = 16'hf6eb;
  rom[32254] = 16'hff2b;
  rom[32255] = 16'hf70a;
  rom[32256] = 16'hff2c;
  rom[32257] = 16'heeab;
  rom[32258] = 16'hff0f;
  rom[32259] = 16'he60c;
  rom[32260] = 16'habc7;
  rom[32261] = 16'h81e2;
  rom[32262] = 16'ha206;
  rom[32263] = 16'hd288;
  rom[32264] = 16'hea29;
  rom[32265] = 16'hf1c7;
  rom[32266] = 16'hf9e7;
  rom[32267] = 16'hf1c6;
  rom[32268] = 16'hea27;
  rom[32269] = 16'hd268;
  rom[32270] = 16'h9a04;
  rom[32271] = 16'h8aa2;
  rom[32272] = 16'hf68c;
  rom[32273] = 16'hfeea;
  rom[32274] = 16'hff6b;
  rom[32275] = 16'hef49;
  rom[32276] = 16'hf729;
  rom[32277] = 16'hf729;
  rom[32278] = 16'hff2a;
  rom[32279] = 16'hff28;
  rom[32280] = 16'hff29;
  rom[32281] = 16'hff28;
  rom[32282] = 16'hff29;
  rom[32283] = 16'hff29;
  rom[32284] = 16'hff29;
  rom[32285] = 16'hff29;
  rom[32286] = 16'hff4a;
  rom[32287] = 16'hff29;
  rom[32288] = 16'hff29;
  rom[32289] = 16'hf729;
  rom[32290] = 16'hff4a;
  rom[32291] = 16'hff29;
  rom[32292] = 16'hff2a;
  rom[32293] = 16'hff28;
  rom[32294] = 16'hff49;
  rom[32295] = 16'hff28;
  rom[32296] = 16'hff08;
  rom[32297] = 16'hff49;
  rom[32298] = 16'hf6e9;
  rom[32299] = 16'hf749;
  rom[32300] = 16'hff6b;
  rom[32301] = 16'hef0d;
  rom[32302] = 16'hacc7;
  rom[32303] = 16'h8363;
  rom[32304] = 16'heead;
  rom[32305] = 16'hf70c;
  rom[32306] = 16'hf729;
  rom[32307] = 16'hf747;
  rom[32308] = 16'hff68;
  rom[32309] = 16'hf709;
  rom[32310] = 16'hff2b;
  rom[32311] = 16'hff0a;
  rom[32312] = 16'hff29;
  rom[32313] = 16'hff28;
  rom[32314] = 16'hff29;
  rom[32315] = 16'hff29;
  rom[32316] = 16'hf72a;
  rom[32317] = 16'hf749;
  rom[32318] = 16'hf74a;
  rom[32319] = 16'hff29;
  rom[32320] = 16'hff2b;
  rom[32321] = 16'hfeca;
  rom[32322] = 16'hff2c;
  rom[32323] = 16'hfeea;
  rom[32324] = 16'hff0c;
  rom[32325] = 16'hc4c8;
  rom[32326] = 16'h8a22;
  rom[32327] = 16'hd287;
  rom[32328] = 16'he246;
  rom[32329] = 16'hd246;
  rom[32330] = 16'hdbad;
  rom[32331] = 16'hff5c;
  rom[32332] = 16'hfffe;
  rom[32333] = 16'hffff;
  rom[32334] = 16'hffff;
  rom[32335] = 16'hffff;
  rom[32336] = 16'hffff;
  rom[32337] = 16'hffff;
  rom[32338] = 16'hffff;
  rom[32339] = 16'hffff;
  rom[32340] = 16'hffff;
  rom[32341] = 16'hffff;
  rom[32342] = 16'hffff;
  rom[32343] = 16'hffff;
  rom[32344] = 16'hffff;
  rom[32345] = 16'hffff;
  rom[32346] = 16'hffff;
  rom[32347] = 16'hffff;
  rom[32348] = 16'hffff;
  rom[32349] = 16'hffff;
  rom[32350] = 16'hffff;
  rom[32351] = 16'hffff;
  rom[32352] = 16'hffff;
  rom[32353] = 16'hffff;
  rom[32354] = 16'hffff;
  rom[32355] = 16'hffff;
  rom[32356] = 16'hffff;
  rom[32357] = 16'hffff;
  rom[32358] = 16'hffff;
  rom[32359] = 16'hffff;
  rom[32360] = 16'hffff;
  rom[32361] = 16'hffff;
  rom[32362] = 16'hffff;
  rom[32363] = 16'hffff;
  rom[32364] = 16'hffff;
  rom[32365] = 16'hffff;
  rom[32366] = 16'hffff;
  rom[32367] = 16'hffff;
  rom[32368] = 16'hffff;
  rom[32369] = 16'hffff;
  rom[32370] = 16'hffff;
  rom[32371] = 16'hffff;
  rom[32372] = 16'hffff;
  rom[32373] = 16'hffff;
  rom[32374] = 16'hffff;
  rom[32375] = 16'hffff;
  rom[32376] = 16'hffff;
  rom[32377] = 16'hffff;
  rom[32378] = 16'hffff;
  rom[32379] = 16'hffff;
  rom[32380] = 16'hffff;
  rom[32381] = 16'hffff;
  rom[32382] = 16'hffff;
  rom[32383] = 16'hffff;
  rom[32384] = 16'hffff;
  rom[32385] = 16'hffff;
  rom[32386] = 16'hffff;
  rom[32387] = 16'hffff;
  rom[32388] = 16'hffff;
  rom[32389] = 16'hffff;
  rom[32390] = 16'hffff;
  rom[32391] = 16'hffff;
  rom[32392] = 16'hffff;
  rom[32393] = 16'hffff;
  rom[32394] = 16'hffff;
  rom[32395] = 16'hffff;
  rom[32396] = 16'hffff;
  rom[32397] = 16'hffff;
  rom[32398] = 16'hffff;
  rom[32399] = 16'hffff;
  rom[32400] = 16'hffff;
  rom[32401] = 16'hffff;
  rom[32402] = 16'hffff;
  rom[32403] = 16'hffff;
  rom[32404] = 16'hffff;
  rom[32405] = 16'hffff;
  rom[32406] = 16'hffff;
  rom[32407] = 16'hffff;
  rom[32408] = 16'hffff;
  rom[32409] = 16'hffff;
  rom[32410] = 16'hffff;
  rom[32411] = 16'hffff;
  rom[32412] = 16'hffff;
  rom[32413] = 16'hffff;
  rom[32414] = 16'hffff;
  rom[32415] = 16'hffff;
  rom[32416] = 16'hffff;
  rom[32417] = 16'hffff;
  rom[32418] = 16'hffff;
  rom[32419] = 16'hffff;
  rom[32420] = 16'hffff;
  rom[32421] = 16'hffff;
  rom[32422] = 16'hffff;
  rom[32423] = 16'hffff;
  rom[32424] = 16'hffde;
  rom[32425] = 16'hffbe;
  rom[32426] = 16'hff5c;
  rom[32427] = 16'hfeda;
  rom[32428] = 16'hed55;
  rom[32429] = 16'hb2eb;
  rom[32430] = 16'hcaeb;
  rom[32431] = 16'hdac9;
  rom[32432] = 16'hca27;
  rom[32433] = 16'he268;
  rom[32434] = 16'hda06;
  rom[32435] = 16'he247;
  rom[32436] = 16'hda26;
  rom[32437] = 16'hd9e5;
  rom[32438] = 16'hd9e5;
  rom[32439] = 16'hea26;
  rom[32440] = 16'hea27;
  rom[32441] = 16'hea06;
  rom[32442] = 16'hd9c5;
  rom[32443] = 16'he1c6;
  rom[32444] = 16'hd9c6;
  rom[32445] = 16'he226;
  rom[32446] = 16'hda46;
  rom[32447] = 16'hca46;
  rom[32448] = 16'hb244;
  rom[32449] = 16'h8141;
  rom[32450] = 16'h58c0;
  rom[32451] = 16'ha324;
  rom[32452] = 16'hf5ee;
  rom[32453] = 16'hfe8f;
  rom[32454] = 16'hf6ae;
  rom[32455] = 16'hfecf;
  rom[32456] = 16'he68e;
  rom[32457] = 16'hde70;
  rom[32458] = 16'h7b44;
  rom[32459] = 16'h59a0;
  rom[32460] = 16'h7203;
  rom[32461] = 16'h9aa7;
  rom[32462] = 16'haa68;
  rom[32463] = 16'hca49;
  rom[32464] = 16'hda28;
  rom[32465] = 16'he9c7;
  rom[32466] = 16'hf206;
  rom[32467] = 16'hf9e6;
  rom[32468] = 16'hf206;
  rom[32469] = 16'he207;
  rom[32470] = 16'hb226;
  rom[32471] = 16'h7a21;
  rom[32472] = 16'hdd69;
  rom[32473] = 16'hfeeb;
  rom[32474] = 16'hf729;
  rom[32475] = 16'hef48;
  rom[32476] = 16'hf708;
  rom[32477] = 16'hff2a;
  rom[32478] = 16'hf709;
  rom[32479] = 16'hf748;
  rom[32480] = 16'hff28;
  rom[32481] = 16'hff48;
  rom[32482] = 16'hf708;
  rom[32483] = 16'hff28;
  rom[32484] = 16'hff08;
  rom[32485] = 16'hff29;
  rom[32486] = 16'hf6e8;
  rom[32487] = 16'hff29;
  rom[32488] = 16'hff29;
  rom[32489] = 16'hff29;
  rom[32490] = 16'hf708;
  rom[32491] = 16'hff29;
  rom[32492] = 16'hff09;
  rom[32493] = 16'hff28;
  rom[32494] = 16'hf728;
  rom[32495] = 16'hff48;
  rom[32496] = 16'hff29;
  rom[32497] = 16'hf6e9;
  rom[32498] = 16'hff8b;
  rom[32499] = 16'hf729;
  rom[32500] = 16'heeea;
  rom[32501] = 16'hd64b;
  rom[32502] = 16'h62a1;
  rom[32503] = 16'hd62c;
  rom[32504] = 16'heeec;
  rom[32505] = 16'hf70a;
  rom[32506] = 16'hf747;
  rom[32507] = 16'hff67;
  rom[32508] = 16'hf747;
  rom[32509] = 16'hff4a;
  rom[32510] = 16'hf70a;
  rom[32511] = 16'hfee9;
  rom[32512] = 16'hfee8;
  rom[32513] = 16'hff28;
  rom[32514] = 16'hf708;
  rom[32515] = 16'hff29;
  rom[32516] = 16'hf729;
  rom[32517] = 16'hf749;
  rom[32518] = 16'hef09;
  rom[32519] = 16'hff29;
  rom[32520] = 16'hfee9;
  rom[32521] = 16'hfeea;
  rom[32522] = 16'hff0a;
  rom[32523] = 16'hf70b;
  rom[32524] = 16'heeec;
  rom[32525] = 16'hc4a8;
  rom[32526] = 16'haa84;
  rom[32527] = 16'hd246;
  rom[32528] = 16'he206;
  rom[32529] = 16'he2a8;
  rom[32530] = 16'hdc4f;
  rom[32531] = 16'hff7c;
  rom[32532] = 16'hffff;
  rom[32533] = 16'hffff;
  rom[32534] = 16'hffdf;
  rom[32535] = 16'hffff;
  rom[32536] = 16'hffff;
  rom[32537] = 16'hffff;
  rom[32538] = 16'hffff;
  rom[32539] = 16'hffff;
  rom[32540] = 16'hffff;
  rom[32541] = 16'hffff;
  rom[32542] = 16'hffff;
  rom[32543] = 16'hffff;
  rom[32544] = 16'hffff;
  rom[32545] = 16'hffff;
  rom[32546] = 16'hffff;
  rom[32547] = 16'hffff;
  rom[32548] = 16'hffff;
  rom[32549] = 16'hffff;
  rom[32550] = 16'hffff;
  rom[32551] = 16'hffff;
  rom[32552] = 16'hffff;
  rom[32553] = 16'hffff;
  rom[32554] = 16'hffff;
  rom[32555] = 16'hffff;
  rom[32556] = 16'hffff;
  rom[32557] = 16'hffff;
  rom[32558] = 16'hffff;
  rom[32559] = 16'hffff;
  rom[32560] = 16'hffff;
  rom[32561] = 16'hffff;
  rom[32562] = 16'hffff;
  rom[32563] = 16'hffff;
  rom[32564] = 16'hffff;
  rom[32565] = 16'hffff;
  rom[32566] = 16'hffff;
  rom[32567] = 16'hffff;
  rom[32568] = 16'hffff;
  rom[32569] = 16'hffff;
  rom[32570] = 16'hffff;
  rom[32571] = 16'hffff;
  rom[32572] = 16'hffff;
  rom[32573] = 16'hffff;
  rom[32574] = 16'hffff;
  rom[32575] = 16'hffff;
  rom[32576] = 16'hffff;
  rom[32577] = 16'hffff;
  rom[32578] = 16'hffff;
  rom[32579] = 16'hffff;
  rom[32580] = 16'hffff;
  rom[32581] = 16'hffff;
  rom[32582] = 16'hffff;
  rom[32583] = 16'hffff;
  rom[32584] = 16'hffff;
  rom[32585] = 16'hffff;
  rom[32586] = 16'hffff;
  rom[32587] = 16'hffff;
  rom[32588] = 16'hffff;
  rom[32589] = 16'hffff;
  rom[32590] = 16'hffff;
  rom[32591] = 16'hffff;
  rom[32592] = 16'hffff;
  rom[32593] = 16'hffff;
  rom[32594] = 16'hffff;
  rom[32595] = 16'hffff;
  rom[32596] = 16'hffff;
  rom[32597] = 16'hffff;
  rom[32598] = 16'hffff;
  rom[32599] = 16'hffff;
  rom[32600] = 16'hffff;
  rom[32601] = 16'hffff;
  rom[32602] = 16'hffff;
  rom[32603] = 16'hffff;
  rom[32604] = 16'hffff;
  rom[32605] = 16'hffff;
  rom[32606] = 16'hffff;
  rom[32607] = 16'hffff;
  rom[32608] = 16'hffff;
  rom[32609] = 16'hffff;
  rom[32610] = 16'hffff;
  rom[32611] = 16'hffff;
  rom[32612] = 16'hffff;
  rom[32613] = 16'hffff;
  rom[32614] = 16'hffff;
  rom[32615] = 16'hffff;
  rom[32616] = 16'hffff;
  rom[32617] = 16'hffff;
  rom[32618] = 16'hffff;
  rom[32619] = 16'hffff;
  rom[32620] = 16'hffff;
  rom[32621] = 16'hffff;
  rom[32622] = 16'hffff;
  rom[32623] = 16'hffff;
  rom[32624] = 16'hffff;
  rom[32625] = 16'hffff;
  rom[32626] = 16'hffff;
  rom[32627] = 16'hff9f;
  rom[32628] = 16'hff7e;
  rom[32629] = 16'hfefc;
  rom[32630] = 16'hedd7;
  rom[32631] = 16'he4d3;
  rom[32632] = 16'hdbef;
  rom[32633] = 16'hcb2b;
  rom[32634] = 16'hd2ea;
  rom[32635] = 16'hd2a9;
  rom[32636] = 16'hdaa9;
  rom[32637] = 16'hda68;
  rom[32638] = 16'hda68;
  rom[32639] = 16'he267;
  rom[32640] = 16'he247;
  rom[32641] = 16'he227;
  rom[32642] = 16'hea68;
  rom[32643] = 16'he227;
  rom[32644] = 16'he228;
  rom[32645] = 16'hda07;
  rom[32646] = 16'he269;
  rom[32647] = 16'hd248;
  rom[32648] = 16'hd2a8;
  rom[32649] = 16'hc2c8;
  rom[32650] = 16'haa86;
  rom[32651] = 16'h8a04;
  rom[32652] = 16'h79e4;
  rom[32653] = 16'h7204;
  rom[32654] = 16'h6a43;
  rom[32655] = 16'h6a43;
  rom[32656] = 16'h6aa6;
  rom[32657] = 16'h72c8;
  rom[32658] = 16'h940c;
  rom[32659] = 16'hb4d0;
  rom[32660] = 16'hcd33;
  rom[32661] = 16'hd512;
  rom[32662] = 16'hd470;
  rom[32663] = 16'hcb8d;
  rom[32664] = 16'hd2eb;
  rom[32665] = 16'hda89;
  rom[32666] = 16'hea48;
  rom[32667] = 16'he9e6;
  rom[32668] = 16'hf227;
  rom[32669] = 16'hea07;
  rom[32670] = 16'hc226;
  rom[32671] = 16'h79a0;
  rom[32672] = 16'hcd08;
  rom[32673] = 16'hff2c;
  rom[32674] = 16'hf768;
  rom[32675] = 16'hef47;
  rom[32676] = 16'hff2a;
  rom[32677] = 16'hfeea;
  rom[32678] = 16'hf72a;
  rom[32679] = 16'hf748;
  rom[32680] = 16'hff49;
  rom[32681] = 16'hf748;
  rom[32682] = 16'hff29;
  rom[32683] = 16'hff28;
  rom[32684] = 16'hff29;
  rom[32685] = 16'hff09;
  rom[32686] = 16'hff2a;
  rom[32687] = 16'hff29;
  rom[32688] = 16'hff29;
  rom[32689] = 16'hff28;
  rom[32690] = 16'hff49;
  rom[32691] = 16'hff29;
  rom[32692] = 16'hff2a;
  rom[32693] = 16'hf729;
  rom[32694] = 16'hff49;
  rom[32695] = 16'hff28;
  rom[32696] = 16'hff2a;
  rom[32697] = 16'hf6e9;
  rom[32698] = 16'hff4a;
  rom[32699] = 16'hef09;
  rom[32700] = 16'hff6d;
  rom[32701] = 16'ha4c6;
  rom[32702] = 16'h9c45;
  rom[32703] = 16'heeed;
  rom[32704] = 16'hf70b;
  rom[32705] = 16'hffeb;
  rom[32706] = 16'hf727;
  rom[32707] = 16'hf727;
  rom[32708] = 16'hff4a;
  rom[32709] = 16'hf72a;
  rom[32710] = 16'hff0a;
  rom[32711] = 16'hff0a;
  rom[32712] = 16'hff2a;
  rom[32713] = 16'hff28;
  rom[32714] = 16'hff48;
  rom[32715] = 16'hf748;
  rom[32716] = 16'hf749;
  rom[32717] = 16'hf729;
  rom[32718] = 16'hff2a;
  rom[32719] = 16'hfee9;
  rom[32720] = 16'hff29;
  rom[32721] = 16'hf708;
  rom[32722] = 16'hf74a;
  rom[32723] = 16'hef2b;
  rom[32724] = 16'he6ad;
  rom[32725] = 16'ha385;
  rom[32726] = 16'hba65;
  rom[32727] = 16'he247;
  rom[32728] = 16'hf227;
  rom[32729] = 16'hd267;
  rom[32730] = 16'hed53;
  rom[32731] = 16'hfffe;
  rom[32732] = 16'hffff;
  rom[32733] = 16'hffff;
  rom[32734] = 16'hffdf;
  rom[32735] = 16'hffff;
  rom[32736] = 16'hffff;
  rom[32737] = 16'hffff;
  rom[32738] = 16'hffff;
  rom[32739] = 16'hffff;
  rom[32740] = 16'hffff;
  rom[32741] = 16'hffff;
  rom[32742] = 16'hffff;
  rom[32743] = 16'hffff;
  rom[32744] = 16'hffff;
  rom[32745] = 16'hffff;
  rom[32746] = 16'hffff;
  rom[32747] = 16'hffff;
  rom[32748] = 16'hffff;
  rom[32749] = 16'hffff;
  rom[32750] = 16'hffff;
  rom[32751] = 16'hffff;
  rom[32752] = 16'hffff;
  rom[32753] = 16'hffff;
  rom[32754] = 16'hffff;
  rom[32755] = 16'hffff;
  rom[32756] = 16'hffff;
  rom[32757] = 16'hffff;
  rom[32758] = 16'hffff;
  rom[32759] = 16'hffff;
  rom[32760] = 16'hffff;
  rom[32761] = 16'hffff;
  rom[32762] = 16'hffff;
  rom[32763] = 16'hffff;
  rom[32764] = 16'hffff;
  rom[32765] = 16'hffff;
  rom[32766] = 16'hffff;
  rom[32767] = 16'hffff;
  rom[32768] = 16'hffff;
  rom[32769] = 16'hffff;
  rom[32770] = 16'hffff;
  rom[32771] = 16'hffff;
  rom[32772] = 16'hffff;
  rom[32773] = 16'hffff;
  rom[32774] = 16'hffff;
  rom[32775] = 16'hffff;
  rom[32776] = 16'hffff;
  rom[32777] = 16'hffff;
  rom[32778] = 16'hffff;
  rom[32779] = 16'hffff;
  rom[32780] = 16'hffff;
  rom[32781] = 16'hffff;
  rom[32782] = 16'hffff;
  rom[32783] = 16'hffff;
  rom[32784] = 16'hffff;
  rom[32785] = 16'hffff;
  rom[32786] = 16'hffff;
  rom[32787] = 16'hffff;
  rom[32788] = 16'hffff;
  rom[32789] = 16'hffff;
  rom[32790] = 16'hffff;
  rom[32791] = 16'hffff;
  rom[32792] = 16'hffff;
  rom[32793] = 16'hffff;
  rom[32794] = 16'hffff;
  rom[32795] = 16'hffff;
  rom[32796] = 16'hffff;
  rom[32797] = 16'hffff;
  rom[32798] = 16'hffff;
  rom[32799] = 16'hffff;
  rom[32800] = 16'hffff;
  rom[32801] = 16'hffff;
  rom[32802] = 16'hffff;
  rom[32803] = 16'hffff;
  rom[32804] = 16'hffff;
  rom[32805] = 16'hffff;
  rom[32806] = 16'hffff;
  rom[32807] = 16'hffff;
  rom[32808] = 16'hffff;
  rom[32809] = 16'hffff;
  rom[32810] = 16'hffff;
  rom[32811] = 16'hffff;
  rom[32812] = 16'hffff;
  rom[32813] = 16'hffff;
  rom[32814] = 16'hffff;
  rom[32815] = 16'hffff;
  rom[32816] = 16'hffff;
  rom[32817] = 16'hffff;
  rom[32818] = 16'hffff;
  rom[32819] = 16'hffff;
  rom[32820] = 16'hffff;
  rom[32821] = 16'hffff;
  rom[32822] = 16'hffff;
  rom[32823] = 16'hffff;
  rom[32824] = 16'hffff;
  rom[32825] = 16'hffff;
  rom[32826] = 16'hffdf;
  rom[32827] = 16'hffff;
  rom[32828] = 16'hffdf;
  rom[32829] = 16'hffbf;
  rom[32830] = 16'hff9e;
  rom[32831] = 16'hff7e;
  rom[32832] = 16'hff1b;
  rom[32833] = 16'hfe99;
  rom[32834] = 16'hfdf7;
  rom[32835] = 16'hf513;
  rom[32836] = 16'hdc30;
  rom[32837] = 16'hd38d;
  rom[32838] = 16'hd32b;
  rom[32839] = 16'hd32b;
  rom[32840] = 16'hd30a;
  rom[32841] = 16'hd30a;
  rom[32842] = 16'hd2ea;
  rom[32843] = 16'hd2ea;
  rom[32844] = 16'hcac9;
  rom[32845] = 16'hdaca;
  rom[32846] = 16'hd2ca;
  rom[32847] = 16'hd30b;
  rom[32848] = 16'hc32a;
  rom[32849] = 16'hc34b;
  rom[32850] = 16'hb36c;
  rom[32851] = 16'hc40e;
  rom[32852] = 16'hc470;
  rom[32853] = 16'hc512;
  rom[32854] = 16'hcdd5;
  rom[32855] = 16'he6b9;
  rom[32856] = 16'hf71b;
  rom[32857] = 16'hff7d;
  rom[32858] = 16'hffbe;
  rom[32859] = 16'hffdf;
  rom[32860] = 16'hffbd;
  rom[32861] = 16'hff9d;
  rom[32862] = 16'hff5b;
  rom[32863] = 16'hfeda;
  rom[32864] = 16'hfdd5;
  rom[32865] = 16'hd3ad;
  rom[32866] = 16'hc248;
  rom[32867] = 16'hda68;
  rom[32868] = 16'hea47;
  rom[32869] = 16'hf1e6;
  rom[32870] = 16'hca06;
  rom[32871] = 16'h8981;
  rom[32872] = 16'hac45;
  rom[32873] = 16'hf70b;
  rom[32874] = 16'hef28;
  rom[32875] = 16'hf748;
  rom[32876] = 16'hfee9;
  rom[32877] = 16'hfeea;
  rom[32878] = 16'hf70a;
  rom[32879] = 16'hf748;
  rom[32880] = 16'hef28;
  rom[32881] = 16'hf748;
  rom[32882] = 16'hff28;
  rom[32883] = 16'hff28;
  rom[32884] = 16'hf708;
  rom[32885] = 16'hff28;
  rom[32886] = 16'hff09;
  rom[32887] = 16'hff29;
  rom[32888] = 16'hf708;
  rom[32889] = 16'hff28;
  rom[32890] = 16'hff08;
  rom[32891] = 16'hff29;
  rom[32892] = 16'hf709;
  rom[32893] = 16'hf729;
  rom[32894] = 16'hf708;
  rom[32895] = 16'hff28;
  rom[32896] = 16'hf709;
  rom[32897] = 16'hff6b;
  rom[32898] = 16'hf70a;
  rom[32899] = 16'hff4c;
  rom[32900] = 16'hd649;
  rom[32901] = 16'h7b61;
  rom[32902] = 16'hd62b;
  rom[32903] = 16'hff4d;
  rom[32904] = 16'hef09;
  rom[32905] = 16'hef07;
  rom[32906] = 16'hf6e7;
  rom[32907] = 16'hff6a;
  rom[32908] = 16'heee8;
  rom[32909] = 16'hff29;
  rom[32910] = 16'hf709;
  rom[32911] = 16'hff0a;
  rom[32912] = 16'hff0a;
  rom[32913] = 16'hff29;
  rom[32914] = 16'hf727;
  rom[32915] = 16'hf747;
  rom[32916] = 16'hf727;
  rom[32917] = 16'hff09;
  rom[32918] = 16'hfee9;
  rom[32919] = 16'hff29;
  rom[32920] = 16'hff27;
  rom[32921] = 16'hf747;
  rom[32922] = 16'hef48;
  rom[32923] = 16'hef2c;
  rom[32924] = 16'hcdcb;
  rom[32925] = 16'h9283;
  rom[32926] = 16'hc225;
  rom[32927] = 16'hfa48;
  rom[32928] = 16'he207;
  rom[32929] = 16'hcaa9;
  rom[32930] = 16'hf637;
  rom[32931] = 16'hfffe;
  rom[32932] = 16'hfffe;
  rom[32933] = 16'hffff;
  rom[32934] = 16'hffbf;
  rom[32935] = 16'hffff;
  rom[32936] = 16'hffff;
  rom[32937] = 16'hffff;
  rom[32938] = 16'hffff;
  rom[32939] = 16'hffff;
  rom[32940] = 16'hffff;
  rom[32941] = 16'hffff;
  rom[32942] = 16'hffff;
  rom[32943] = 16'hffff;
  rom[32944] = 16'hffff;
  rom[32945] = 16'hffff;
  rom[32946] = 16'hffff;
  rom[32947] = 16'hffff;
  rom[32948] = 16'hffff;
  rom[32949] = 16'hffff;
  rom[32950] = 16'hffff;
  rom[32951] = 16'hffff;
  rom[32952] = 16'hffff;
  rom[32953] = 16'hffff;
  rom[32954] = 16'hffff;
  rom[32955] = 16'hffff;
  rom[32956] = 16'hffff;
  rom[32957] = 16'hffff;
  rom[32958] = 16'hffff;
  rom[32959] = 16'hffff;
  rom[32960] = 16'hffff;
  rom[32961] = 16'hffff;
  rom[32962] = 16'hffff;
  rom[32963] = 16'hffff;
  rom[32964] = 16'hffff;
  rom[32965] = 16'hffff;
  rom[32966] = 16'hffff;
  rom[32967] = 16'hffff;
  rom[32968] = 16'hffff;
  rom[32969] = 16'hffff;
  rom[32970] = 16'hffff;
  rom[32971] = 16'hffff;
  rom[32972] = 16'hffff;
  rom[32973] = 16'hffff;
  rom[32974] = 16'hffff;
  rom[32975] = 16'hffff;
  rom[32976] = 16'hffff;
  rom[32977] = 16'hffff;
  rom[32978] = 16'hffff;
  rom[32979] = 16'hffff;
  rom[32980] = 16'hffff;
  rom[32981] = 16'hffff;
  rom[32982] = 16'hffff;
  rom[32983] = 16'hffff;
  rom[32984] = 16'hffff;
  rom[32985] = 16'hffff;
  rom[32986] = 16'hffff;
  rom[32987] = 16'hffff;
  rom[32988] = 16'hffff;
  rom[32989] = 16'hffff;
  rom[32990] = 16'hffff;
  rom[32991] = 16'hffff;
  rom[32992] = 16'hffff;
  rom[32993] = 16'hffff;
  rom[32994] = 16'hffff;
  rom[32995] = 16'hffff;
  rom[32996] = 16'hffff;
  rom[32997] = 16'hffff;
  rom[32998] = 16'hffff;
  rom[32999] = 16'hffff;
  rom[33000] = 16'hffff;
  rom[33001] = 16'hffff;
  rom[33002] = 16'hffff;
  rom[33003] = 16'hffff;
  rom[33004] = 16'hffff;
  rom[33005] = 16'hffff;
  rom[33006] = 16'hffff;
  rom[33007] = 16'hffff;
  rom[33008] = 16'hffff;
  rom[33009] = 16'hffff;
  rom[33010] = 16'hffff;
  rom[33011] = 16'hffff;
  rom[33012] = 16'hffff;
  rom[33013] = 16'hffff;
  rom[33014] = 16'hffff;
  rom[33015] = 16'hffff;
  rom[33016] = 16'hffff;
  rom[33017] = 16'hffff;
  rom[33018] = 16'hffff;
  rom[33019] = 16'hffff;
  rom[33020] = 16'hffff;
  rom[33021] = 16'hffff;
  rom[33022] = 16'hffff;
  rom[33023] = 16'hffff;
  rom[33024] = 16'hffff;
  rom[33025] = 16'hffff;
  rom[33026] = 16'hffff;
  rom[33027] = 16'hffff;
  rom[33028] = 16'hffff;
  rom[33029] = 16'hffff;
  rom[33030] = 16'hffff;
  rom[33031] = 16'hffff;
  rom[33032] = 16'hffff;
  rom[33033] = 16'hffdf;
  rom[33034] = 16'hffff;
  rom[33035] = 16'hff7d;
  rom[33036] = 16'hff7d;
  rom[33037] = 16'hff3c;
  rom[33038] = 16'hff3c;
  rom[33039] = 16'hfe99;
  rom[33040] = 16'hfe58;
  rom[33041] = 16'hf617;
  rom[33042] = 16'hf637;
  rom[33043] = 16'hf616;
  rom[33044] = 16'hf637;
  rom[33045] = 16'hf636;
  rom[33046] = 16'hf616;
  rom[33047] = 16'hf637;
  rom[33048] = 16'hfe98;
  rom[33049] = 16'hfeb9;
  rom[33050] = 16'hff5c;
  rom[33051] = 16'hff9d;
  rom[33052] = 16'hffdf;
  rom[33053] = 16'hffbe;
  rom[33054] = 16'hffff;
  rom[33055] = 16'hffff;
  rom[33056] = 16'hffff;
  rom[33057] = 16'hffff;
  rom[33058] = 16'hffff;
  rom[33059] = 16'hffdf;
  rom[33060] = 16'hffff;
  rom[33061] = 16'hffdf;
  rom[33062] = 16'hffff;
  rom[33063] = 16'hffde;
  rom[33064] = 16'hffbe;
  rom[33065] = 16'hff1b;
  rom[33066] = 16'hf575;
  rom[33067] = 16'hcb2b;
  rom[33068] = 16'hda88;
  rom[33069] = 16'he228;
  rom[33070] = 16'hda68;
  rom[33071] = 16'h99c2;
  rom[33072] = 16'h9343;
  rom[33073] = 16'he6ab;
  rom[33074] = 16'he729;
  rom[33075] = 16'hff28;
  rom[33076] = 16'hfee9;
  rom[33077] = 16'hfeea;
  rom[33078] = 16'hff2a;
  rom[33079] = 16'hf748;
  rom[33080] = 16'hf749;
  rom[33081] = 16'hf748;
  rom[33082] = 16'hff29;
  rom[33083] = 16'hff28;
  rom[33084] = 16'hff29;
  rom[33085] = 16'hff28;
  rom[33086] = 16'hff29;
  rom[33087] = 16'hff28;
  rom[33088] = 16'hff29;
  rom[33089] = 16'hff28;
  rom[33090] = 16'hff29;
  rom[33091] = 16'hff29;
  rom[33092] = 16'hff2a;
  rom[33093] = 16'hf729;
  rom[33094] = 16'hff2a;
  rom[33095] = 16'hff29;
  rom[33096] = 16'hff09;
  rom[33097] = 16'hff0a;
  rom[33098] = 16'hf6ea;
  rom[33099] = 16'hf74d;
  rom[33100] = 16'ha4c5;
  rom[33101] = 16'h9c65;
  rom[33102] = 16'hf6ed;
  rom[33103] = 16'hef0a;
  rom[33104] = 16'hff69;
  rom[33105] = 16'hf748;
  rom[33106] = 16'hf74a;
  rom[33107] = 16'hff4b;
  rom[33108] = 16'hf70a;
  rom[33109] = 16'hf729;
  rom[33110] = 16'hff29;
  rom[33111] = 16'hff09;
  rom[33112] = 16'hff2a;
  rom[33113] = 16'hf729;
  rom[33114] = 16'hf748;
  rom[33115] = 16'hf747;
  rom[33116] = 16'hff28;
  rom[33117] = 16'hff09;
  rom[33118] = 16'hff0a;
  rom[33119] = 16'hff09;
  rom[33120] = 16'hff47;
  rom[33121] = 16'hf747;
  rom[33122] = 16'hf76a;
  rom[33123] = 16'hf72d;
  rom[33124] = 16'hc4ea;
  rom[33125] = 16'ha284;
  rom[33126] = 16'he288;
  rom[33127] = 16'he9c7;
  rom[33128] = 16'hea69;
  rom[33129] = 16'hd36c;
  rom[33130] = 16'hff3b;
  rom[33131] = 16'hffde;
  rom[33132] = 16'hffff;
  rom[33133] = 16'hffff;
  rom[33134] = 16'hffff;
  rom[33135] = 16'hffff;
  rom[33136] = 16'hffff;
  rom[33137] = 16'hffff;
  rom[33138] = 16'hffff;
  rom[33139] = 16'hffff;
  rom[33140] = 16'hffff;
  rom[33141] = 16'hffff;
  rom[33142] = 16'hffff;
  rom[33143] = 16'hffff;
  rom[33144] = 16'hffff;
  rom[33145] = 16'hffff;
  rom[33146] = 16'hffff;
  rom[33147] = 16'hffff;
  rom[33148] = 16'hffff;
  rom[33149] = 16'hffff;
  rom[33150] = 16'hffff;
  rom[33151] = 16'hffff;
  rom[33152] = 16'hffff;
  rom[33153] = 16'hffff;
  rom[33154] = 16'hffff;
  rom[33155] = 16'hffff;
  rom[33156] = 16'hffff;
  rom[33157] = 16'hffff;
  rom[33158] = 16'hffff;
  rom[33159] = 16'hffff;
  rom[33160] = 16'hffff;
  rom[33161] = 16'hffff;
  rom[33162] = 16'hffff;
  rom[33163] = 16'hffff;
  rom[33164] = 16'hffff;
  rom[33165] = 16'hffff;
  rom[33166] = 16'hffff;
  rom[33167] = 16'hffff;
  rom[33168] = 16'hffff;
  rom[33169] = 16'hffff;
  rom[33170] = 16'hffff;
  rom[33171] = 16'hffff;
  rom[33172] = 16'hffff;
  rom[33173] = 16'hffff;
  rom[33174] = 16'hffff;
  rom[33175] = 16'hffff;
  rom[33176] = 16'hffff;
  rom[33177] = 16'hffff;
  rom[33178] = 16'hffff;
  rom[33179] = 16'hffff;
  rom[33180] = 16'hffff;
  rom[33181] = 16'hffff;
  rom[33182] = 16'hffff;
  rom[33183] = 16'hffff;
  rom[33184] = 16'hffff;
  rom[33185] = 16'hffff;
  rom[33186] = 16'hffff;
  rom[33187] = 16'hffff;
  rom[33188] = 16'hffff;
  rom[33189] = 16'hffff;
  rom[33190] = 16'hffff;
  rom[33191] = 16'hffff;
  rom[33192] = 16'hffff;
  rom[33193] = 16'hffff;
  rom[33194] = 16'hffff;
  rom[33195] = 16'hffff;
  rom[33196] = 16'hffff;
  rom[33197] = 16'hffff;
  rom[33198] = 16'hffff;
  rom[33199] = 16'hffff;
  rom[33200] = 16'hffff;
  rom[33201] = 16'hffff;
  rom[33202] = 16'hffff;
  rom[33203] = 16'hffff;
  rom[33204] = 16'hffff;
  rom[33205] = 16'hffff;
  rom[33206] = 16'hffff;
  rom[33207] = 16'hffff;
  rom[33208] = 16'hffff;
  rom[33209] = 16'hffff;
  rom[33210] = 16'hffff;
  rom[33211] = 16'hffff;
  rom[33212] = 16'hffff;
  rom[33213] = 16'hffff;
  rom[33214] = 16'hffff;
  rom[33215] = 16'hffff;
  rom[33216] = 16'hffff;
  rom[33217] = 16'hffff;
  rom[33218] = 16'hffff;
  rom[33219] = 16'hffff;
  rom[33220] = 16'hffff;
  rom[33221] = 16'hffff;
  rom[33222] = 16'hffff;
  rom[33223] = 16'hffff;
  rom[33224] = 16'hffff;
  rom[33225] = 16'hffff;
  rom[33226] = 16'hfffe;
  rom[33227] = 16'hffff;
  rom[33228] = 16'hffff;
  rom[33229] = 16'hffff;
  rom[33230] = 16'hffff;
  rom[33231] = 16'hffff;
  rom[33232] = 16'hffff;
  rom[33233] = 16'hffff;
  rom[33234] = 16'hffff;
  rom[33235] = 16'hffff;
  rom[33236] = 16'hffdf;
  rom[33237] = 16'hffdf;
  rom[33238] = 16'hffdf;
  rom[33239] = 16'hffdf;
  rom[33240] = 16'hffbe;
  rom[33241] = 16'hffdf;
  rom[33242] = 16'hffde;
  rom[33243] = 16'hffde;
  rom[33244] = 16'hffbe;
  rom[33245] = 16'hfffe;
  rom[33246] = 16'hfffd;
  rom[33247] = 16'hfffe;
  rom[33248] = 16'hffde;
  rom[33249] = 16'hffff;
  rom[33250] = 16'hffdf;
  rom[33251] = 16'hffff;
  rom[33252] = 16'hffdf;
  rom[33253] = 16'hffff;
  rom[33254] = 16'hffff;
  rom[33255] = 16'hffff;
  rom[33256] = 16'hffde;
  rom[33257] = 16'hfffe;
  rom[33258] = 16'hffff;
  rom[33259] = 16'hffff;
  rom[33260] = 16'hffff;
  rom[33261] = 16'hffff;
  rom[33262] = 16'hffff;
  rom[33263] = 16'hffdf;
  rom[33264] = 16'hffbe;
  rom[33265] = 16'hffdf;
  rom[33266] = 16'hff5c;
  rom[33267] = 16'hfe37;
  rom[33268] = 16'hdbce;
  rom[33269] = 16'hd28a;
  rom[33270] = 16'hca47;
  rom[33271] = 16'ha204;
  rom[33272] = 16'h7a22;
  rom[33273] = 16'he68c;
  rom[33274] = 16'he729;
  rom[33275] = 16'hff29;
  rom[33276] = 16'hfec9;
  rom[33277] = 16'hff0a;
  rom[33278] = 16'hf709;
  rom[33279] = 16'hf748;
  rom[33280] = 16'hf728;
  rom[33281] = 16'hf748;
  rom[33282] = 16'hf708;
  rom[33283] = 16'hff29;
  rom[33284] = 16'hff09;
  rom[33285] = 16'hff29;
  rom[33286] = 16'hf708;
  rom[33287] = 16'hff28;
  rom[33288] = 16'hff08;
  rom[33289] = 16'hff28;
  rom[33290] = 16'hf708;
  rom[33291] = 16'hff29;
  rom[33292] = 16'hff09;
  rom[33293] = 16'hff29;
  rom[33294] = 16'hf709;
  rom[33295] = 16'hff29;
  rom[33296] = 16'hff29;
  rom[33297] = 16'hff2a;
  rom[33298] = 16'hf70a;
  rom[33299] = 16'heecc;
  rom[33300] = 16'h7b60;
  rom[33301] = 16'hbd47;
  rom[33302] = 16'hef0b;
  rom[33303] = 16'hf72a;
  rom[33304] = 16'hf727;
  rom[33305] = 16'hff48;
  rom[33306] = 16'hf708;
  rom[33307] = 16'hf72b;
  rom[33308] = 16'hf70a;
  rom[33309] = 16'hf72a;
  rom[33310] = 16'hf708;
  rom[33311] = 16'hff49;
  rom[33312] = 16'hff09;
  rom[33313] = 16'hff29;
  rom[33314] = 16'hef27;
  rom[33315] = 16'hff47;
  rom[33316] = 16'hff08;
  rom[33317] = 16'hff0a;
  rom[33318] = 16'hff0a;
  rom[33319] = 16'hf708;
  rom[33320] = 16'hf748;
  rom[33321] = 16'hf728;
  rom[33322] = 16'heeea;
  rom[33323] = 16'hee2c;
  rom[33324] = 16'h8aa3;
  rom[33325] = 16'hb246;
  rom[33326] = 16'hd206;
  rom[33327] = 16'he248;
  rom[33328] = 16'hc248;
  rom[33329] = 16'hecf2;
  rom[33330] = 16'hff9d;
  rom[33331] = 16'hffff;
  rom[33332] = 16'hffff;
  rom[33333] = 16'hffff;
  rom[33334] = 16'hffdf;
  rom[33335] = 16'hffff;
  rom[33336] = 16'hffff;
  rom[33337] = 16'hffff;
  rom[33338] = 16'hffff;
  rom[33339] = 16'hffff;
  rom[33340] = 16'hffff;
  rom[33341] = 16'hffff;
  rom[33342] = 16'hffff;
  rom[33343] = 16'hffff;
  rom[33344] = 16'hffff;
  rom[33345] = 16'hffff;
  rom[33346] = 16'hffff;
  rom[33347] = 16'hffff;
  rom[33348] = 16'hffff;
  rom[33349] = 16'hffff;
  rom[33350] = 16'hffff;
  rom[33351] = 16'hffff;
  rom[33352] = 16'hffff;
  rom[33353] = 16'hffff;
  rom[33354] = 16'hffff;
  rom[33355] = 16'hffff;
  rom[33356] = 16'hffff;
  rom[33357] = 16'hffff;
  rom[33358] = 16'hffff;
  rom[33359] = 16'hffff;
  rom[33360] = 16'hffff;
  rom[33361] = 16'hffff;
  rom[33362] = 16'hffff;
  rom[33363] = 16'hffff;
  rom[33364] = 16'hffff;
  rom[33365] = 16'hffff;
  rom[33366] = 16'hffff;
  rom[33367] = 16'hffff;
  rom[33368] = 16'hffff;
  rom[33369] = 16'hffff;
  rom[33370] = 16'hffff;
  rom[33371] = 16'hffff;
  rom[33372] = 16'hffff;
  rom[33373] = 16'hffff;
  rom[33374] = 16'hffff;
  rom[33375] = 16'hffff;
  rom[33376] = 16'hffff;
  rom[33377] = 16'hffff;
  rom[33378] = 16'hffff;
  rom[33379] = 16'hffff;
  rom[33380] = 16'hffff;
  rom[33381] = 16'hffff;
  rom[33382] = 16'hffff;
  rom[33383] = 16'hffff;
  rom[33384] = 16'hffff;
  rom[33385] = 16'hffff;
  rom[33386] = 16'hffff;
  rom[33387] = 16'hffff;
  rom[33388] = 16'hffff;
  rom[33389] = 16'hffff;
  rom[33390] = 16'hffff;
  rom[33391] = 16'hffff;
  rom[33392] = 16'hffff;
  rom[33393] = 16'hffff;
  rom[33394] = 16'hffff;
  rom[33395] = 16'hffff;
  rom[33396] = 16'hffff;
  rom[33397] = 16'hffff;
  rom[33398] = 16'hffff;
  rom[33399] = 16'hffff;
  rom[33400] = 16'hffff;
  rom[33401] = 16'hffff;
  rom[33402] = 16'hffff;
  rom[33403] = 16'hffff;
  rom[33404] = 16'hffff;
  rom[33405] = 16'hffff;
  rom[33406] = 16'hffff;
  rom[33407] = 16'hffff;
  rom[33408] = 16'hffff;
  rom[33409] = 16'hffff;
  rom[33410] = 16'hffff;
  rom[33411] = 16'hffff;
  rom[33412] = 16'hffff;
  rom[33413] = 16'hffff;
  rom[33414] = 16'hffff;
  rom[33415] = 16'hffff;
  rom[33416] = 16'hffff;
  rom[33417] = 16'hffff;
  rom[33418] = 16'hffff;
  rom[33419] = 16'hffff;
  rom[33420] = 16'hffff;
  rom[33421] = 16'hffff;
  rom[33422] = 16'hffff;
  rom[33423] = 16'hffff;
  rom[33424] = 16'hffff;
  rom[33425] = 16'hffff;
  rom[33426] = 16'hffff;
  rom[33427] = 16'hffff;
  rom[33428] = 16'hffdf;
  rom[33429] = 16'hffff;
  rom[33430] = 16'hffff;
  rom[33431] = 16'hffff;
  rom[33432] = 16'hffff;
  rom[33433] = 16'hffff;
  rom[33434] = 16'hffdf;
  rom[33435] = 16'hffff;
  rom[33436] = 16'hffff;
  rom[33437] = 16'hffff;
  rom[33438] = 16'hffdf;
  rom[33439] = 16'hffdf;
  rom[33440] = 16'hffff;
  rom[33441] = 16'hffff;
  rom[33442] = 16'hffff;
  rom[33443] = 16'hffff;
  rom[33444] = 16'hffff;
  rom[33445] = 16'hffff;
  rom[33446] = 16'hffff;
  rom[33447] = 16'hffff;
  rom[33448] = 16'hffff;
  rom[33449] = 16'hffff;
  rom[33450] = 16'hffff;
  rom[33451] = 16'hffff;
  rom[33452] = 16'hffff;
  rom[33453] = 16'hffdf;
  rom[33454] = 16'hffff;
  rom[33455] = 16'hffdf;
  rom[33456] = 16'hffff;
  rom[33457] = 16'hffdf;
  rom[33458] = 16'hffff;
  rom[33459] = 16'hffff;
  rom[33460] = 16'hffff;
  rom[33461] = 16'hffff;
  rom[33462] = 16'hffdf;
  rom[33463] = 16'hffbf;
  rom[33464] = 16'hffff;
  rom[33465] = 16'hffff;
  rom[33466] = 16'hffdf;
  rom[33467] = 16'hff9e;
  rom[33468] = 16'hfe59;
  rom[33469] = 16'hcb6e;
  rom[33470] = 16'hcaeb;
  rom[33471] = 16'ha205;
  rom[33472] = 16'h79e2;
  rom[33473] = 16'hd5eb;
  rom[33474] = 16'hf74c;
  rom[33475] = 16'hf709;
  rom[33476] = 16'hff0a;
  rom[33477] = 16'hff09;
  rom[33478] = 16'hff49;
  rom[33479] = 16'hf748;
  rom[33480] = 16'hf749;
  rom[33481] = 16'hf748;
  rom[33482] = 16'hff29;
  rom[33483] = 16'hff29;
  rom[33484] = 16'hff2a;
  rom[33485] = 16'hff29;
  rom[33486] = 16'hff29;
  rom[33487] = 16'hff28;
  rom[33488] = 16'hff29;
  rom[33489] = 16'hff28;
  rom[33490] = 16'hff29;
  rom[33491] = 16'hff29;
  rom[33492] = 16'hff29;
  rom[33493] = 16'hff29;
  rom[33494] = 16'hff2a;
  rom[33495] = 16'hff29;
  rom[33496] = 16'hff29;
  rom[33497] = 16'hf709;
  rom[33498] = 16'hff2c;
  rom[33499] = 16'hc587;
  rom[33500] = 16'h8be2;
  rom[33501] = 16'hd62a;
  rom[33502] = 16'hff2d;
  rom[33503] = 16'hf729;
  rom[33504] = 16'hf729;
  rom[33505] = 16'hff28;
  rom[33506] = 16'hff49;
  rom[33507] = 16'hff29;
  rom[33508] = 16'hf70a;
  rom[33509] = 16'hff49;
  rom[33510] = 16'hff49;
  rom[33511] = 16'hf729;
  rom[33512] = 16'hff4a;
  rom[33513] = 16'hf728;
  rom[33514] = 16'hf749;
  rom[33515] = 16'hff27;
  rom[33516] = 16'hff29;
  rom[33517] = 16'hff0a;
  rom[33518] = 16'hff0a;
  rom[33519] = 16'hff49;
  rom[33520] = 16'hf749;
  rom[33521] = 16'hff4a;
  rom[33522] = 16'hfeac;
  rom[33523] = 16'hc447;
  rom[33524] = 16'h9a24;
  rom[33525] = 16'hca47;
  rom[33526] = 16'hea68;
  rom[33527] = 16'hda47;
  rom[33528] = 16'hcb0b;
  rom[33529] = 16'hf657;
  rom[33530] = 16'hffde;
  rom[33531] = 16'hffff;
  rom[33532] = 16'hffff;
  rom[33533] = 16'hffff;
  rom[33534] = 16'hffff;
  rom[33535] = 16'hffff;
  rom[33536] = 16'hffff;
  rom[33537] = 16'hffff;
  rom[33538] = 16'hffff;
  rom[33539] = 16'hffff;
  rom[33540] = 16'hffff;
  rom[33541] = 16'hffff;
  rom[33542] = 16'hffff;
  rom[33543] = 16'hffff;
  rom[33544] = 16'hffff;
  rom[33545] = 16'hffff;
  rom[33546] = 16'hffff;
  rom[33547] = 16'hffff;
  rom[33548] = 16'hffff;
  rom[33549] = 16'hffff;
  rom[33550] = 16'hffff;
  rom[33551] = 16'hffff;
  rom[33552] = 16'hffff;
  rom[33553] = 16'hffff;
  rom[33554] = 16'hffff;
  rom[33555] = 16'hffff;
  rom[33556] = 16'hffff;
  rom[33557] = 16'hffff;
  rom[33558] = 16'hffff;
  rom[33559] = 16'hffff;
  rom[33560] = 16'hffff;
  rom[33561] = 16'hffff;
  rom[33562] = 16'hffff;
  rom[33563] = 16'hffff;
  rom[33564] = 16'hffff;
  rom[33565] = 16'hffff;
  rom[33566] = 16'hffff;
  rom[33567] = 16'hffff;
  rom[33568] = 16'hffff;
  rom[33569] = 16'hffff;
  rom[33570] = 16'hffff;
  rom[33571] = 16'hffff;
  rom[33572] = 16'hffff;
  rom[33573] = 16'hffff;
  rom[33574] = 16'hffff;
  rom[33575] = 16'hffff;
  rom[33576] = 16'hffff;
  rom[33577] = 16'hffff;
  rom[33578] = 16'hffff;
  rom[33579] = 16'hffff;
  rom[33580] = 16'hffff;
  rom[33581] = 16'hffff;
  rom[33582] = 16'hffff;
  rom[33583] = 16'hffff;
  rom[33584] = 16'hffff;
  rom[33585] = 16'hffff;
  rom[33586] = 16'hffff;
  rom[33587] = 16'hffff;
  rom[33588] = 16'hffff;
  rom[33589] = 16'hffff;
  rom[33590] = 16'hffff;
  rom[33591] = 16'hffff;
  rom[33592] = 16'hffff;
  rom[33593] = 16'hffff;
  rom[33594] = 16'hffff;
  rom[33595] = 16'hffff;
  rom[33596] = 16'hffff;
  rom[33597] = 16'hffff;
  rom[33598] = 16'hffff;
  rom[33599] = 16'hffff;
  rom[33600] = 16'hffff;
  rom[33601] = 16'hffff;
  rom[33602] = 16'hffff;
  rom[33603] = 16'hffff;
  rom[33604] = 16'hffff;
  rom[33605] = 16'hffff;
  rom[33606] = 16'hffff;
  rom[33607] = 16'hffff;
  rom[33608] = 16'hffff;
  rom[33609] = 16'hffff;
  rom[33610] = 16'hffff;
  rom[33611] = 16'hffff;
  rom[33612] = 16'hffff;
  rom[33613] = 16'hffff;
  rom[33614] = 16'hffff;
  rom[33615] = 16'hffff;
  rom[33616] = 16'hffff;
  rom[33617] = 16'hffff;
  rom[33618] = 16'hffff;
  rom[33619] = 16'hffff;
  rom[33620] = 16'hffff;
  rom[33621] = 16'hffff;
  rom[33622] = 16'hffff;
  rom[33623] = 16'hffff;
  rom[33624] = 16'hffff;
  rom[33625] = 16'hffff;
  rom[33626] = 16'hffff;
  rom[33627] = 16'hffff;
  rom[33628] = 16'hffdf;
  rom[33629] = 16'hffff;
  rom[33630] = 16'hf7ff;
  rom[33631] = 16'hffff;
  rom[33632] = 16'hffff;
  rom[33633] = 16'hffff;
  rom[33634] = 16'hffff;
  rom[33635] = 16'hffff;
  rom[33636] = 16'hffff;
  rom[33637] = 16'hffff;
  rom[33638] = 16'hffff;
  rom[33639] = 16'hffff;
  rom[33640] = 16'hffff;
  rom[33641] = 16'hffff;
  rom[33642] = 16'hffff;
  rom[33643] = 16'hffff;
  rom[33644] = 16'hffff;
  rom[33645] = 16'hffff;
  rom[33646] = 16'hffff;
  rom[33647] = 16'hffff;
  rom[33648] = 16'hffff;
  rom[33649] = 16'hffff;
  rom[33650] = 16'hffff;
  rom[33651] = 16'hffff;
  rom[33652] = 16'hffff;
  rom[33653] = 16'hffff;
  rom[33654] = 16'hffdf;
  rom[33655] = 16'hffdf;
  rom[33656] = 16'hffdf;
  rom[33657] = 16'hffff;
  rom[33658] = 16'hf7ff;
  rom[33659] = 16'hffff;
  rom[33660] = 16'hffff;
  rom[33661] = 16'hffff;
  rom[33662] = 16'hffff;
  rom[33663] = 16'hffff;
  rom[33664] = 16'hffdf;
  rom[33665] = 16'hffff;
  rom[33666] = 16'hffff;
  rom[33667] = 16'hffbf;
  rom[33668] = 16'hff7e;
  rom[33669] = 16'hfe7a;
  rom[33670] = 16'hd3ef;
  rom[33671] = 16'hbaca;
  rom[33672] = 16'h79a1;
  rom[33673] = 16'hbca8;
  rom[33674] = 16'hf72c;
  rom[33675] = 16'hf72a;
  rom[33676] = 16'hf709;
  rom[33677] = 16'hff09;
  rom[33678] = 16'hff29;
  rom[33679] = 16'hff28;
  rom[33680] = 16'hf728;
  rom[33681] = 16'hf728;
  rom[33682] = 16'hff09;
  rom[33683] = 16'hff29;
  rom[33684] = 16'hf709;
  rom[33685] = 16'hff29;
  rom[33686] = 16'hff08;
  rom[33687] = 16'hff28;
  rom[33688] = 16'hf708;
  rom[33689] = 16'hff28;
  rom[33690] = 16'hff08;
  rom[33691] = 16'hff28;
  rom[33692] = 16'hf728;
  rom[33693] = 16'hff29;
  rom[33694] = 16'hff09;
  rom[33695] = 16'hff2a;
  rom[33696] = 16'hf729;
  rom[33697] = 16'hf709;
  rom[33698] = 16'hf70b;
  rom[33699] = 16'hacc5;
  rom[33700] = 16'h9c43;
  rom[33701] = 16'heeec;
  rom[33702] = 16'hef0b;
  rom[33703] = 16'hff2a;
  rom[33704] = 16'hf729;
  rom[33705] = 16'hff49;
  rom[33706] = 16'hf708;
  rom[33707] = 16'hff29;
  rom[33708] = 16'hf729;
  rom[33709] = 16'hf729;
  rom[33710] = 16'hf728;
  rom[33711] = 16'hff29;
  rom[33712] = 16'hf708;
  rom[33713] = 16'hff48;
  rom[33714] = 16'hff28;
  rom[33715] = 16'hff29;
  rom[33716] = 16'hf709;
  rom[33717] = 16'hff0a;
  rom[33718] = 16'hf709;
  rom[33719] = 16'hff2a;
  rom[33720] = 16'hef09;
  rom[33721] = 16'hf6ec;
  rom[33722] = 16'hedeb;
  rom[33723] = 16'ha2a3;
  rom[33724] = 16'hb225;
  rom[33725] = 16'he288;
  rom[33726] = 16'hda06;
  rom[33727] = 16'hd289;
  rom[33728] = 16'hdc70;
  rom[33729] = 16'hff7c;
  rom[33730] = 16'hffdf;
  rom[33731] = 16'hffff;
  rom[33732] = 16'hffdf;
  rom[33733] = 16'hffff;
  rom[33734] = 16'hffff;
  rom[33735] = 16'hffff;
  rom[33736] = 16'hffff;
  rom[33737] = 16'hffff;
  rom[33738] = 16'hffff;
  rom[33739] = 16'hffff;
  rom[33740] = 16'hffff;
  rom[33741] = 16'hffff;
  rom[33742] = 16'hffff;
  rom[33743] = 16'hffff;
  rom[33744] = 16'hffff;
  rom[33745] = 16'hffff;
  rom[33746] = 16'hffff;
  rom[33747] = 16'hffff;
  rom[33748] = 16'hffff;
  rom[33749] = 16'hffff;
  rom[33750] = 16'hffff;
  rom[33751] = 16'hffff;
  rom[33752] = 16'hffff;
  rom[33753] = 16'hffff;
  rom[33754] = 16'hffff;
  rom[33755] = 16'hffff;
  rom[33756] = 16'hffff;
  rom[33757] = 16'hffff;
  rom[33758] = 16'hffff;
  rom[33759] = 16'hffff;
  rom[33760] = 16'hffff;
  rom[33761] = 16'hffff;
  rom[33762] = 16'hffff;
  rom[33763] = 16'hffff;
  rom[33764] = 16'hffff;
  rom[33765] = 16'hffff;
  rom[33766] = 16'hffff;
  rom[33767] = 16'hffff;
  rom[33768] = 16'hffff;
  rom[33769] = 16'hffff;
  rom[33770] = 16'hffff;
  rom[33771] = 16'hffff;
  rom[33772] = 16'hffff;
  rom[33773] = 16'hffff;
  rom[33774] = 16'hffff;
  rom[33775] = 16'hffff;
  rom[33776] = 16'hffff;
  rom[33777] = 16'hffff;
  rom[33778] = 16'hffff;
  rom[33779] = 16'hffff;
  rom[33780] = 16'hffff;
  rom[33781] = 16'hffff;
  rom[33782] = 16'hffff;
  rom[33783] = 16'hffff;
  rom[33784] = 16'hffff;
  rom[33785] = 16'hffff;
  rom[33786] = 16'hffff;
  rom[33787] = 16'hffff;
  rom[33788] = 16'hffff;
  rom[33789] = 16'hffff;
  rom[33790] = 16'hffff;
  rom[33791] = 16'hffff;
  rom[33792] = 16'hffff;
  rom[33793] = 16'hffff;
  rom[33794] = 16'hffff;
  rom[33795] = 16'hffff;
  rom[33796] = 16'hffff;
  rom[33797] = 16'hffff;
  rom[33798] = 16'hffff;
  rom[33799] = 16'hffff;
  rom[33800] = 16'hffff;
  rom[33801] = 16'hffff;
  rom[33802] = 16'hffff;
  rom[33803] = 16'hffff;
  rom[33804] = 16'hffff;
  rom[33805] = 16'hffff;
  rom[33806] = 16'hffff;
  rom[33807] = 16'hffff;
  rom[33808] = 16'hffff;
  rom[33809] = 16'hffff;
  rom[33810] = 16'hffff;
  rom[33811] = 16'hffff;
  rom[33812] = 16'hffff;
  rom[33813] = 16'hffff;
  rom[33814] = 16'hffff;
  rom[33815] = 16'hffff;
  rom[33816] = 16'hffff;
  rom[33817] = 16'hffff;
  rom[33818] = 16'hffff;
  rom[33819] = 16'hffff;
  rom[33820] = 16'hffff;
  rom[33821] = 16'hffff;
  rom[33822] = 16'hffff;
  rom[33823] = 16'hffff;
  rom[33824] = 16'hffff;
  rom[33825] = 16'hffff;
  rom[33826] = 16'hffff;
  rom[33827] = 16'hffff;
  rom[33828] = 16'hffff;
  rom[33829] = 16'hffff;
  rom[33830] = 16'hffff;
  rom[33831] = 16'hffff;
  rom[33832] = 16'hffff;
  rom[33833] = 16'hffff;
  rom[33834] = 16'hffff;
  rom[33835] = 16'hffff;
  rom[33836] = 16'hffff;
  rom[33837] = 16'hffff;
  rom[33838] = 16'hffff;
  rom[33839] = 16'hffff;
  rom[33840] = 16'hffff;
  rom[33841] = 16'hffff;
  rom[33842] = 16'hffff;
  rom[33843] = 16'hffff;
  rom[33844] = 16'hffff;
  rom[33845] = 16'hffff;
  rom[33846] = 16'hffff;
  rom[33847] = 16'hffff;
  rom[33848] = 16'hffff;
  rom[33849] = 16'hffff;
  rom[33850] = 16'hffff;
  rom[33851] = 16'hffff;
  rom[33852] = 16'hffff;
  rom[33853] = 16'hffff;
  rom[33854] = 16'hffff;
  rom[33855] = 16'hffff;
  rom[33856] = 16'hffff;
  rom[33857] = 16'hffff;
  rom[33858] = 16'hffff;
  rom[33859] = 16'hffff;
  rom[33860] = 16'hffff;
  rom[33861] = 16'hffff;
  rom[33862] = 16'hffff;
  rom[33863] = 16'hffff;
  rom[33864] = 16'hffff;
  rom[33865] = 16'hffff;
  rom[33866] = 16'hffff;
  rom[33867] = 16'hffff;
  rom[33868] = 16'hffdf;
  rom[33869] = 16'hff9d;
  rom[33870] = 16'hfdf7;
  rom[33871] = 16'hc38d;
  rom[33872] = 16'h7183;
  rom[33873] = 16'hac07;
  rom[33874] = 16'hf6ed;
  rom[33875] = 16'hf74b;
  rom[33876] = 16'hf74a;
  rom[33877] = 16'hff29;
  rom[33878] = 16'hff09;
  rom[33879] = 16'hff28;
  rom[33880] = 16'hff29;
  rom[33881] = 16'hff29;
  rom[33882] = 16'hff2a;
  rom[33883] = 16'hff29;
  rom[33884] = 16'hff2a;
  rom[33885] = 16'hff29;
  rom[33886] = 16'hff2a;
  rom[33887] = 16'hff29;
  rom[33888] = 16'hff29;
  rom[33889] = 16'hff28;
  rom[33890] = 16'hff49;
  rom[33891] = 16'hf747;
  rom[33892] = 16'hff29;
  rom[33893] = 16'hff29;
  rom[33894] = 16'hff0b;
  rom[33895] = 16'hff0a;
  rom[33896] = 16'hff29;
  rom[33897] = 16'hf709;
  rom[33898] = 16'hf70c;
  rom[33899] = 16'h9c64;
  rom[33900] = 16'hbd67;
  rom[33901] = 16'hf72b;
  rom[33902] = 16'hef2a;
  rom[33903] = 16'hf729;
  rom[33904] = 16'hf72a;
  rom[33905] = 16'hff49;
  rom[33906] = 16'hff29;
  rom[33907] = 16'hff28;
  rom[33908] = 16'hff29;
  rom[33909] = 16'hff28;
  rom[33910] = 16'hff29;
  rom[33911] = 16'hff28;
  rom[33912] = 16'hff29;
  rom[33913] = 16'hef28;
  rom[33914] = 16'hf749;
  rom[33915] = 16'hff2a;
  rom[33916] = 16'hff0a;
  rom[33917] = 16'hff29;
  rom[33918] = 16'hff49;
  rom[33919] = 16'hf728;
  rom[33920] = 16'hff4c;
  rom[33921] = 16'hf66c;
  rom[33922] = 16'hdcea;
  rom[33923] = 16'h9a03;
  rom[33924] = 16'hd2a6;
  rom[33925] = 16'hea87;
  rom[33926] = 16'hda07;
  rom[33927] = 16'hd32b;
  rom[33928] = 16'hfe38;
  rom[33929] = 16'hff9d;
  rom[33930] = 16'hffff;
  rom[33931] = 16'hffff;
  rom[33932] = 16'hffff;
  rom[33933] = 16'hffff;
  rom[33934] = 16'hffff;
  rom[33935] = 16'hffff;
  rom[33936] = 16'hffff;
  rom[33937] = 16'hffff;
  rom[33938] = 16'hffff;
  rom[33939] = 16'hffff;
  rom[33940] = 16'hffff;
  rom[33941] = 16'hffff;
  rom[33942] = 16'hffff;
  rom[33943] = 16'hffff;
  rom[33944] = 16'hffff;
  rom[33945] = 16'hffff;
  rom[33946] = 16'hffff;
  rom[33947] = 16'hffff;
  rom[33948] = 16'hffff;
  rom[33949] = 16'hffff;
  rom[33950] = 16'hffff;
  rom[33951] = 16'hffff;
  rom[33952] = 16'hffff;
  rom[33953] = 16'hffff;
  rom[33954] = 16'hffff;
  rom[33955] = 16'hffff;
  rom[33956] = 16'hffff;
  rom[33957] = 16'hffff;
  rom[33958] = 16'hffff;
  rom[33959] = 16'hffff;
  rom[33960] = 16'hffff;
  rom[33961] = 16'hffff;
  rom[33962] = 16'hffff;
  rom[33963] = 16'hffff;
  rom[33964] = 16'hffff;
  rom[33965] = 16'hffff;
  rom[33966] = 16'hffff;
  rom[33967] = 16'hffff;
  rom[33968] = 16'hffff;
  rom[33969] = 16'hffff;
  rom[33970] = 16'hffff;
  rom[33971] = 16'hffff;
  rom[33972] = 16'hffff;
  rom[33973] = 16'hffff;
  rom[33974] = 16'hffff;
  rom[33975] = 16'hffff;
  rom[33976] = 16'hffff;
  rom[33977] = 16'hffff;
  rom[33978] = 16'hffff;
  rom[33979] = 16'hffff;
  rom[33980] = 16'hffff;
  rom[33981] = 16'hffff;
  rom[33982] = 16'hffff;
  rom[33983] = 16'hffff;
  rom[33984] = 16'hffff;
  rom[33985] = 16'hffff;
  rom[33986] = 16'hffff;
  rom[33987] = 16'hffff;
  rom[33988] = 16'hffff;
  rom[33989] = 16'hffff;
  rom[33990] = 16'hffff;
  rom[33991] = 16'hffff;
  rom[33992] = 16'hffff;
  rom[33993] = 16'hffff;
  rom[33994] = 16'hffff;
  rom[33995] = 16'hffff;
  rom[33996] = 16'hffff;
  rom[33997] = 16'hffff;
  rom[33998] = 16'hffff;
  rom[33999] = 16'hffff;
  rom[34000] = 16'hffff;
  rom[34001] = 16'hffff;
  rom[34002] = 16'hffff;
  rom[34003] = 16'hffff;
  rom[34004] = 16'hffff;
  rom[34005] = 16'hffff;
  rom[34006] = 16'hffff;
  rom[34007] = 16'hffff;
  rom[34008] = 16'hffff;
  rom[34009] = 16'hffff;
  rom[34010] = 16'hffff;
  rom[34011] = 16'hffff;
  rom[34012] = 16'hffff;
  rom[34013] = 16'hffff;
  rom[34014] = 16'hffff;
  rom[34015] = 16'hffff;
  rom[34016] = 16'hffff;
  rom[34017] = 16'hffff;
  rom[34018] = 16'hffff;
  rom[34019] = 16'hffff;
  rom[34020] = 16'hffff;
  rom[34021] = 16'hffff;
  rom[34022] = 16'hffff;
  rom[34023] = 16'hffff;
  rom[34024] = 16'hffff;
  rom[34025] = 16'hffff;
  rom[34026] = 16'hffff;
  rom[34027] = 16'hffff;
  rom[34028] = 16'hffff;
  rom[34029] = 16'hffff;
  rom[34030] = 16'hffff;
  rom[34031] = 16'hffff;
  rom[34032] = 16'hffff;
  rom[34033] = 16'hffff;
  rom[34034] = 16'hffff;
  rom[34035] = 16'hffff;
  rom[34036] = 16'hffff;
  rom[34037] = 16'hffff;
  rom[34038] = 16'hffff;
  rom[34039] = 16'hffff;
  rom[34040] = 16'hffff;
  rom[34041] = 16'hffff;
  rom[34042] = 16'hffff;
  rom[34043] = 16'hffff;
  rom[34044] = 16'hffff;
  rom[34045] = 16'hffff;
  rom[34046] = 16'hffff;
  rom[34047] = 16'hffff;
  rom[34048] = 16'hffff;
  rom[34049] = 16'hffff;
  rom[34050] = 16'hffff;
  rom[34051] = 16'hffff;
  rom[34052] = 16'hffff;
  rom[34053] = 16'hffff;
  rom[34054] = 16'hffff;
  rom[34055] = 16'hffff;
  rom[34056] = 16'hffff;
  rom[34057] = 16'hffff;
  rom[34058] = 16'hffff;
  rom[34059] = 16'hffff;
  rom[34060] = 16'hffff;
  rom[34061] = 16'hffff;
  rom[34062] = 16'hffdf;
  rom[34063] = 16'hffff;
  rom[34064] = 16'hffff;
  rom[34065] = 16'hffff;
  rom[34066] = 16'hffff;
  rom[34067] = 16'hffff;
  rom[34068] = 16'hffff;
  rom[34069] = 16'hffbe;
  rom[34070] = 16'hfefb;
  rom[34071] = 16'hdd14;
  rom[34072] = 16'h8266;
  rom[34073] = 16'h9345;
  rom[34074] = 16'heecd;
  rom[34075] = 16'hf70a;
  rom[34076] = 16'hef29;
  rom[34077] = 16'hff29;
  rom[34078] = 16'hff08;
  rom[34079] = 16'hff28;
  rom[34080] = 16'hff08;
  rom[34081] = 16'hff29;
  rom[34082] = 16'hf708;
  rom[34083] = 16'hff29;
  rom[34084] = 16'hff09;
  rom[34085] = 16'hff29;
  rom[34086] = 16'hf709;
  rom[34087] = 16'hff29;
  rom[34088] = 16'hff08;
  rom[34089] = 16'hff28;
  rom[34090] = 16'hf727;
  rom[34091] = 16'hf748;
  rom[34092] = 16'hff28;
  rom[34093] = 16'hff29;
  rom[34094] = 16'hf6ea;
  rom[34095] = 16'hff0a;
  rom[34096] = 16'hf708;
  rom[34097] = 16'hf729;
  rom[34098] = 16'he6ab;
  rom[34099] = 16'ha485;
  rom[34100] = 16'hce0a;
  rom[34101] = 16'hf72c;
  rom[34102] = 16'hf74a;
  rom[34103] = 16'hf749;
  rom[34104] = 16'hf729;
  rom[34105] = 16'hff29;
  rom[34106] = 16'hf729;
  rom[34107] = 16'hff29;
  rom[34108] = 16'hff08;
  rom[34109] = 16'hff29;
  rom[34110] = 16'hf708;
  rom[34111] = 16'hff29;
  rom[34112] = 16'hff08;
  rom[34113] = 16'hff49;
  rom[34114] = 16'hf728;
  rom[34115] = 16'hf729;
  rom[34116] = 16'hf729;
  rom[34117] = 16'hf728;
  rom[34118] = 16'hf728;
  rom[34119] = 16'hef2a;
  rom[34120] = 16'hf6ed;
  rom[34121] = 16'he58c;
  rom[34122] = 16'h9a83;
  rom[34123] = 16'hba86;
  rom[34124] = 16'hda86;
  rom[34125] = 16'hda46;
  rom[34126] = 16'hd2a8;
  rom[34127] = 16'hecb1;
  rom[34128] = 16'hff1b;
  rom[34129] = 16'hffff;
  rom[34130] = 16'hffdf;
  rom[34131] = 16'hffff;
  rom[34132] = 16'hffff;
  rom[34133] = 16'hffff;
  rom[34134] = 16'hffff;
  rom[34135] = 16'hffff;
  rom[34136] = 16'hffff;
  rom[34137] = 16'hffff;
  rom[34138] = 16'hffff;
  rom[34139] = 16'hffff;
  rom[34140] = 16'hffff;
  rom[34141] = 16'hffff;
  rom[34142] = 16'hffff;
  rom[34143] = 16'hffff;
  rom[34144] = 16'hffff;
  rom[34145] = 16'hffff;
  rom[34146] = 16'hffff;
  rom[34147] = 16'hffff;
  rom[34148] = 16'hffff;
  rom[34149] = 16'hffff;
  rom[34150] = 16'hffff;
  rom[34151] = 16'hffff;
  rom[34152] = 16'hffff;
  rom[34153] = 16'hffff;
  rom[34154] = 16'hffff;
  rom[34155] = 16'hffff;
  rom[34156] = 16'hffff;
  rom[34157] = 16'hffff;
  rom[34158] = 16'hffff;
  rom[34159] = 16'hffff;
  rom[34160] = 16'hffff;
  rom[34161] = 16'hffff;
  rom[34162] = 16'hffff;
  rom[34163] = 16'hffff;
  rom[34164] = 16'hffff;
  rom[34165] = 16'hffff;
  rom[34166] = 16'hffff;
  rom[34167] = 16'hffff;
  rom[34168] = 16'hffff;
  rom[34169] = 16'hffff;
  rom[34170] = 16'hffff;
  rom[34171] = 16'hffff;
  rom[34172] = 16'hffff;
  rom[34173] = 16'hffff;
  rom[34174] = 16'hffff;
  rom[34175] = 16'hffff;
  rom[34176] = 16'hffff;
  rom[34177] = 16'hffff;
  rom[34178] = 16'hffff;
  rom[34179] = 16'hffff;
  rom[34180] = 16'hffff;
  rom[34181] = 16'hffff;
  rom[34182] = 16'hffff;
  rom[34183] = 16'hffff;
  rom[34184] = 16'hffff;
  rom[34185] = 16'hffff;
  rom[34186] = 16'hffff;
  rom[34187] = 16'hffff;
  rom[34188] = 16'hffff;
  rom[34189] = 16'hffff;
  rom[34190] = 16'hffff;
  rom[34191] = 16'hffff;
  rom[34192] = 16'hffff;
  rom[34193] = 16'hffff;
  rom[34194] = 16'hffff;
  rom[34195] = 16'hffff;
  rom[34196] = 16'hffff;
  rom[34197] = 16'hffff;
  rom[34198] = 16'hffff;
  rom[34199] = 16'hffff;
  rom[34200] = 16'hffff;
  rom[34201] = 16'hffff;
  rom[34202] = 16'hffff;
  rom[34203] = 16'hffff;
  rom[34204] = 16'hffff;
  rom[34205] = 16'hffff;
  rom[34206] = 16'hffff;
  rom[34207] = 16'hffff;
  rom[34208] = 16'hffff;
  rom[34209] = 16'hffff;
  rom[34210] = 16'hffff;
  rom[34211] = 16'hffff;
  rom[34212] = 16'hffff;
  rom[34213] = 16'hffff;
  rom[34214] = 16'hffff;
  rom[34215] = 16'hffff;
  rom[34216] = 16'hffff;
  rom[34217] = 16'hffff;
  rom[34218] = 16'hffff;
  rom[34219] = 16'hffff;
  rom[34220] = 16'hffff;
  rom[34221] = 16'hffff;
  rom[34222] = 16'hffff;
  rom[34223] = 16'hffff;
  rom[34224] = 16'hffff;
  rom[34225] = 16'hffff;
  rom[34226] = 16'hffff;
  rom[34227] = 16'hffff;
  rom[34228] = 16'hffff;
  rom[34229] = 16'hffff;
  rom[34230] = 16'hffff;
  rom[34231] = 16'hffff;
  rom[34232] = 16'hffff;
  rom[34233] = 16'hffff;
  rom[34234] = 16'hffff;
  rom[34235] = 16'hffff;
  rom[34236] = 16'hffff;
  rom[34237] = 16'hffff;
  rom[34238] = 16'hffff;
  rom[34239] = 16'hffff;
  rom[34240] = 16'hffff;
  rom[34241] = 16'hffff;
  rom[34242] = 16'hffff;
  rom[34243] = 16'hffff;
  rom[34244] = 16'hffff;
  rom[34245] = 16'hffff;
  rom[34246] = 16'hffff;
  rom[34247] = 16'hffff;
  rom[34248] = 16'hffff;
  rom[34249] = 16'hffff;
  rom[34250] = 16'hffff;
  rom[34251] = 16'hffff;
  rom[34252] = 16'hffff;
  rom[34253] = 16'hffff;
  rom[34254] = 16'hffff;
  rom[34255] = 16'hffff;
  rom[34256] = 16'hffff;
  rom[34257] = 16'hffff;
  rom[34258] = 16'hffff;
  rom[34259] = 16'hffff;
  rom[34260] = 16'hffff;
  rom[34261] = 16'hffff;
  rom[34262] = 16'hffff;
  rom[34263] = 16'hffff;
  rom[34264] = 16'hffff;
  rom[34265] = 16'hffff;
  rom[34266] = 16'hffff;
  rom[34267] = 16'hffff;
  rom[34268] = 16'hffff;
  rom[34269] = 16'hffff;
  rom[34270] = 16'hffdf;
  rom[34271] = 16'hfefb;
  rom[34272] = 16'hb44f;
  rom[34273] = 16'h6a62;
  rom[34274] = 16'he64c;
  rom[34275] = 16'hf70b;
  rom[34276] = 16'hf70a;
  rom[34277] = 16'hff2a;
  rom[34278] = 16'hff09;
  rom[34279] = 16'hff28;
  rom[34280] = 16'hff29;
  rom[34281] = 16'hff28;
  rom[34282] = 16'hff29;
  rom[34283] = 16'hff29;
  rom[34284] = 16'hff2a;
  rom[34285] = 16'hff29;
  rom[34286] = 16'hff2a;
  rom[34287] = 16'hff29;
  rom[34288] = 16'hff29;
  rom[34289] = 16'hff28;
  rom[34290] = 16'hff29;
  rom[34291] = 16'hff28;
  rom[34292] = 16'hff29;
  rom[34293] = 16'hff28;
  rom[34294] = 16'hff2a;
  rom[34295] = 16'hff0a;
  rom[34296] = 16'hff29;
  rom[34297] = 16'hf709;
  rom[34298] = 16'heecb;
  rom[34299] = 16'h9403;
  rom[34300] = 16'hde4b;
  rom[34301] = 16'hf72c;
  rom[34302] = 16'hff6a;
  rom[34303] = 16'hf729;
  rom[34304] = 16'hff4a;
  rom[34305] = 16'hf729;
  rom[34306] = 16'hff4a;
  rom[34307] = 16'hff29;
  rom[34308] = 16'hff29;
  rom[34309] = 16'hff28;
  rom[34310] = 16'hff2a;
  rom[34311] = 16'hf729;
  rom[34312] = 16'hff2a;
  rom[34313] = 16'hff29;
  rom[34314] = 16'hff29;
  rom[34315] = 16'hff49;
  rom[34316] = 16'hff69;
  rom[34317] = 16'hff6a;
  rom[34318] = 16'hf72a;
  rom[34319] = 16'hff2d;
  rom[34320] = 16'he64d;
  rom[34321] = 16'h9b24;
  rom[34322] = 16'h91e3;
  rom[34323] = 16'hc287;
  rom[34324] = 16'hd226;
  rom[34325] = 16'hd288;
  rom[34326] = 16'he42e;
  rom[34327] = 16'hfe78;
  rom[34328] = 16'hffdd;
  rom[34329] = 16'hffff;
  rom[34330] = 16'hffff;
  rom[34331] = 16'hffff;
  rom[34332] = 16'hffff;
  rom[34333] = 16'hffff;
  rom[34334] = 16'hffff;
  rom[34335] = 16'hffff;
  rom[34336] = 16'hffff;
  rom[34337] = 16'hffff;
  rom[34338] = 16'hffff;
  rom[34339] = 16'hffff;
  rom[34340] = 16'hffff;
  rom[34341] = 16'hffff;
  rom[34342] = 16'hffff;
  rom[34343] = 16'hffff;
  rom[34344] = 16'hffff;
  rom[34345] = 16'hffff;
  rom[34346] = 16'hffff;
  rom[34347] = 16'hffff;
  rom[34348] = 16'hffff;
  rom[34349] = 16'hffff;
  rom[34350] = 16'hffff;
  rom[34351] = 16'hffff;
  rom[34352] = 16'hffff;
  rom[34353] = 16'hffff;
  rom[34354] = 16'hffff;
  rom[34355] = 16'hffff;
  rom[34356] = 16'hffff;
  rom[34357] = 16'hffff;
  rom[34358] = 16'hffff;
  rom[34359] = 16'hffff;
  rom[34360] = 16'hffff;
  rom[34361] = 16'hffff;
  rom[34362] = 16'hffff;
  rom[34363] = 16'hffff;
  rom[34364] = 16'hffff;
  rom[34365] = 16'hffff;
  rom[34366] = 16'hffff;
  rom[34367] = 16'hffff;
  rom[34368] = 16'hffff;
  rom[34369] = 16'hffff;
  rom[34370] = 16'hffff;
  rom[34371] = 16'hffff;
  rom[34372] = 16'hffff;
  rom[34373] = 16'hffff;
  rom[34374] = 16'hffff;
  rom[34375] = 16'hffff;
  rom[34376] = 16'hffff;
  rom[34377] = 16'hffff;
  rom[34378] = 16'hffff;
  rom[34379] = 16'hffff;
  rom[34380] = 16'hffff;
  rom[34381] = 16'hffff;
  rom[34382] = 16'hffff;
  rom[34383] = 16'hffff;
  rom[34384] = 16'hffff;
  rom[34385] = 16'hffff;
  rom[34386] = 16'hffff;
  rom[34387] = 16'hffff;
  rom[34388] = 16'hffff;
  rom[34389] = 16'hffff;
  rom[34390] = 16'hffff;
  rom[34391] = 16'hffff;
  rom[34392] = 16'hffff;
  rom[34393] = 16'hffff;
  rom[34394] = 16'hffff;
  rom[34395] = 16'hffff;
  rom[34396] = 16'hffff;
  rom[34397] = 16'hffff;
  rom[34398] = 16'hffff;
  rom[34399] = 16'hffff;
  rom[34400] = 16'hffff;
  rom[34401] = 16'hffff;
  rom[34402] = 16'hffff;
  rom[34403] = 16'hffff;
  rom[34404] = 16'hffff;
  rom[34405] = 16'hffff;
  rom[34406] = 16'hffff;
  rom[34407] = 16'hffff;
  rom[34408] = 16'hffff;
  rom[34409] = 16'hffff;
  rom[34410] = 16'hffff;
  rom[34411] = 16'hffff;
  rom[34412] = 16'hffff;
  rom[34413] = 16'hffff;
  rom[34414] = 16'hffff;
  rom[34415] = 16'hffff;
  rom[34416] = 16'hffff;
  rom[34417] = 16'hffff;
  rom[34418] = 16'hffff;
  rom[34419] = 16'hffff;
  rom[34420] = 16'hffff;
  rom[34421] = 16'hffff;
  rom[34422] = 16'hffff;
  rom[34423] = 16'hffff;
  rom[34424] = 16'hffff;
  rom[34425] = 16'hffff;
  rom[34426] = 16'hffff;
  rom[34427] = 16'hffff;
  rom[34428] = 16'hffff;
  rom[34429] = 16'hffff;
  rom[34430] = 16'hffff;
  rom[34431] = 16'hffff;
  rom[34432] = 16'hffff;
  rom[34433] = 16'hffff;
  rom[34434] = 16'hffff;
  rom[34435] = 16'hffff;
  rom[34436] = 16'hffff;
  rom[34437] = 16'hffff;
  rom[34438] = 16'hffff;
  rom[34439] = 16'hffff;
  rom[34440] = 16'hffff;
  rom[34441] = 16'hffff;
  rom[34442] = 16'hffff;
  rom[34443] = 16'hffff;
  rom[34444] = 16'hffff;
  rom[34445] = 16'hffff;
  rom[34446] = 16'hffff;
  rom[34447] = 16'hffff;
  rom[34448] = 16'hffff;
  rom[34449] = 16'hffff;
  rom[34450] = 16'hffff;
  rom[34451] = 16'hffff;
  rom[34452] = 16'hffff;
  rom[34453] = 16'hffff;
  rom[34454] = 16'hffff;
  rom[34455] = 16'hffff;
  rom[34456] = 16'hffff;
  rom[34457] = 16'hffff;
  rom[34458] = 16'hffff;
  rom[34459] = 16'hffff;
  rom[34460] = 16'hffff;
  rom[34461] = 16'hffff;
  rom[34462] = 16'hffff;
  rom[34463] = 16'hffff;
  rom[34464] = 16'hffff;
  rom[34465] = 16'hffff;
  rom[34466] = 16'hffff;
  rom[34467] = 16'hffff;
  rom[34468] = 16'hffff;
  rom[34469] = 16'hffff;
  rom[34470] = 16'hffdf;
  rom[34471] = 16'hffff;
  rom[34472] = 16'hcdf5;
  rom[34473] = 16'h62a4;
  rom[34474] = 16'hc58a;
  rom[34475] = 16'hfeec;
  rom[34476] = 16'hf70a;
  rom[34477] = 16'hff2a;
  rom[34478] = 16'hf72a;
  rom[34479] = 16'hff28;
  rom[34480] = 16'hf708;
  rom[34481] = 16'hff28;
  rom[34482] = 16'hff08;
  rom[34483] = 16'hff28;
  rom[34484] = 16'hf708;
  rom[34485] = 16'hff28;
  rom[34486] = 16'hff08;
  rom[34487] = 16'hff28;
  rom[34488] = 16'hf708;
  rom[34489] = 16'hff28;
  rom[34490] = 16'hff08;
  rom[34491] = 16'hff29;
  rom[34492] = 16'hf709;
  rom[34493] = 16'hff28;
  rom[34494] = 16'hff08;
  rom[34495] = 16'hff09;
  rom[34496] = 16'hf708;
  rom[34497] = 16'hf729;
  rom[34498] = 16'he6ab;
  rom[34499] = 16'h8ba3;
  rom[34500] = 16'hde4b;
  rom[34501] = 16'hff4c;
  rom[34502] = 16'hf74a;
  rom[34503] = 16'hf729;
  rom[34504] = 16'hf729;
  rom[34505] = 16'hf728;
  rom[34506] = 16'hff28;
  rom[34507] = 16'hff28;
  rom[34508] = 16'hf708;
  rom[34509] = 16'hff28;
  rom[34510] = 16'hf728;
  rom[34511] = 16'hf748;
  rom[34512] = 16'hf708;
  rom[34513] = 16'hfee9;
  rom[34514] = 16'hf708;
  rom[34515] = 16'hf727;
  rom[34516] = 16'hef48;
  rom[34517] = 16'he709;
  rom[34518] = 16'hf72d;
  rom[34519] = 16'hfeef;
  rom[34520] = 16'hb427;
  rom[34521] = 16'h91e2;
  rom[34522] = 16'hcae8;
  rom[34523] = 16'hda68;
  rom[34524] = 16'hdaa9;
  rom[34525] = 16'hd34c;
  rom[34526] = 16'hfe16;
  rom[34527] = 16'hff7c;
  rom[34528] = 16'hffdd;
  rom[34529] = 16'hffff;
  rom[34530] = 16'hffff;
  rom[34531] = 16'hffff;
  rom[34532] = 16'hffff;
  rom[34533] = 16'hffff;
  rom[34534] = 16'hffff;
  rom[34535] = 16'hffff;
  rom[34536] = 16'hffff;
  rom[34537] = 16'hffff;
  rom[34538] = 16'hffff;
  rom[34539] = 16'hffff;
  rom[34540] = 16'hffff;
  rom[34541] = 16'hffff;
  rom[34542] = 16'hffff;
  rom[34543] = 16'hffff;
  rom[34544] = 16'hffff;
  rom[34545] = 16'hffff;
  rom[34546] = 16'hffff;
  rom[34547] = 16'hffff;
  rom[34548] = 16'hffff;
  rom[34549] = 16'hffff;
  rom[34550] = 16'hffff;
  rom[34551] = 16'hffff;
  rom[34552] = 16'hffff;
  rom[34553] = 16'hffff;
  rom[34554] = 16'hffff;
  rom[34555] = 16'hffff;
  rom[34556] = 16'hffff;
  rom[34557] = 16'hffff;
  rom[34558] = 16'hffff;
  rom[34559] = 16'hffff;
  rom[34560] = 16'hffff;
  rom[34561] = 16'hffff;
  rom[34562] = 16'hffff;
  rom[34563] = 16'hffff;
  rom[34564] = 16'hffff;
  rom[34565] = 16'hffff;
  rom[34566] = 16'hffff;
  rom[34567] = 16'hffff;
  rom[34568] = 16'hffff;
  rom[34569] = 16'hffff;
  rom[34570] = 16'hffff;
  rom[34571] = 16'hffff;
  rom[34572] = 16'hffff;
  rom[34573] = 16'hffff;
  rom[34574] = 16'hffff;
  rom[34575] = 16'hffff;
  rom[34576] = 16'hffff;
  rom[34577] = 16'hffff;
  rom[34578] = 16'hffff;
  rom[34579] = 16'hffff;
  rom[34580] = 16'hffff;
  rom[34581] = 16'hffff;
  rom[34582] = 16'hffff;
  rom[34583] = 16'hffff;
  rom[34584] = 16'hffff;
  rom[34585] = 16'hffff;
  rom[34586] = 16'hffff;
  rom[34587] = 16'hffff;
  rom[34588] = 16'hffff;
  rom[34589] = 16'hffff;
  rom[34590] = 16'hffff;
  rom[34591] = 16'hffff;
  rom[34592] = 16'hffff;
  rom[34593] = 16'hffff;
  rom[34594] = 16'hffff;
  rom[34595] = 16'hffff;
  rom[34596] = 16'hffff;
  rom[34597] = 16'hffff;
  rom[34598] = 16'hffff;
  rom[34599] = 16'hffff;
  rom[34600] = 16'hffff;
  rom[34601] = 16'hffff;
  rom[34602] = 16'hffff;
  rom[34603] = 16'hffff;
  rom[34604] = 16'hffff;
  rom[34605] = 16'hffff;
  rom[34606] = 16'hffff;
  rom[34607] = 16'hffff;
  rom[34608] = 16'hffff;
  rom[34609] = 16'hffff;
  rom[34610] = 16'hffff;
  rom[34611] = 16'hffff;
  rom[34612] = 16'hffff;
  rom[34613] = 16'hffff;
  rom[34614] = 16'hffff;
  rom[34615] = 16'hffff;
  rom[34616] = 16'hffff;
  rom[34617] = 16'hffff;
  rom[34618] = 16'hffff;
  rom[34619] = 16'hffff;
  rom[34620] = 16'hffff;
  rom[34621] = 16'hffff;
  rom[34622] = 16'hffff;
  rom[34623] = 16'hffff;
  rom[34624] = 16'hffff;
  rom[34625] = 16'hffff;
  rom[34626] = 16'hffff;
  rom[34627] = 16'hffff;
  rom[34628] = 16'hffff;
  rom[34629] = 16'hffff;
  rom[34630] = 16'hffff;
  rom[34631] = 16'hffff;
  rom[34632] = 16'hffff;
  rom[34633] = 16'hffff;
  rom[34634] = 16'hffff;
  rom[34635] = 16'hffff;
  rom[34636] = 16'hffff;
  rom[34637] = 16'hffff;
  rom[34638] = 16'hffff;
  rom[34639] = 16'hffff;
  rom[34640] = 16'hffff;
  rom[34641] = 16'hffff;
  rom[34642] = 16'hffff;
  rom[34643] = 16'hffff;
  rom[34644] = 16'hffff;
  rom[34645] = 16'hffff;
  rom[34646] = 16'hffff;
  rom[34647] = 16'hffff;
  rom[34648] = 16'hffff;
  rom[34649] = 16'hffff;
  rom[34650] = 16'hffff;
  rom[34651] = 16'hffff;
  rom[34652] = 16'hffff;
  rom[34653] = 16'hffff;
  rom[34654] = 16'hffff;
  rom[34655] = 16'hffff;
  rom[34656] = 16'hffff;
  rom[34657] = 16'hffff;
  rom[34658] = 16'hffff;
  rom[34659] = 16'hffff;
  rom[34660] = 16'hffff;
  rom[34661] = 16'hffff;
  rom[34662] = 16'hffff;
  rom[34663] = 16'hffff;
  rom[34664] = 16'hffff;
  rom[34665] = 16'hffff;
  rom[34666] = 16'hffff;
  rom[34667] = 16'hffff;
  rom[34668] = 16'hffff;
  rom[34669] = 16'hffff;
  rom[34670] = 16'hffff;
  rom[34671] = 16'hffff;
  rom[34672] = 16'hef3b;
  rom[34673] = 16'h7327;
  rom[34674] = 16'hb4c9;
  rom[34675] = 16'hfeed;
  rom[34676] = 16'hff0b;
  rom[34677] = 16'hf709;
  rom[34678] = 16'hff2a;
  rom[34679] = 16'hff28;
  rom[34680] = 16'hff29;
  rom[34681] = 16'hff28;
  rom[34682] = 16'hff29;
  rom[34683] = 16'hff28;
  rom[34684] = 16'hff29;
  rom[34685] = 16'hff28;
  rom[34686] = 16'hff29;
  rom[34687] = 16'hff28;
  rom[34688] = 16'hff29;
  rom[34689] = 16'hff28;
  rom[34690] = 16'hff29;
  rom[34691] = 16'hff29;
  rom[34692] = 16'hff2a;
  rom[34693] = 16'hff27;
  rom[34694] = 16'hff29;
  rom[34695] = 16'hff09;
  rom[34696] = 16'hff2a;
  rom[34697] = 16'hf72a;
  rom[34698] = 16'he68b;
  rom[34699] = 16'h8bc3;
  rom[34700] = 16'he6ad;
  rom[34701] = 16'hf72b;
  rom[34702] = 16'hff6a;
  rom[34703] = 16'hf729;
  rom[34704] = 16'hff29;
  rom[34705] = 16'hf728;
  rom[34706] = 16'hff29;
  rom[34707] = 16'hff28;
  rom[34708] = 16'hff29;
  rom[34709] = 16'hff28;
  rom[34710] = 16'hff29;
  rom[34711] = 16'hf728;
  rom[34712] = 16'hff29;
  rom[34713] = 16'hff0a;
  rom[34714] = 16'hff4a;
  rom[34715] = 16'hf708;
  rom[34716] = 16'hf78b;
  rom[34717] = 16'hdf2b;
  rom[34718] = 16'hf72f;
  rom[34719] = 16'hbc89;
  rom[34720] = 16'h9223;
  rom[34721] = 16'hc2a6;
  rom[34722] = 16'hda88;
  rom[34723] = 16'hd268;
  rom[34724] = 16'hd2aa;
  rom[34725] = 16'hf595;
  rom[34726] = 16'hff5b;
  rom[34727] = 16'hfffe;
  rom[34728] = 16'hffff;
  rom[34729] = 16'hffff;
  rom[34730] = 16'hffff;
  rom[34731] = 16'hffff;
  rom[34732] = 16'hffff;
  rom[34733] = 16'hffff;
  rom[34734] = 16'hffff;
  rom[34735] = 16'hffff;
  rom[34736] = 16'hffff;
  rom[34737] = 16'hffff;
  rom[34738] = 16'hffff;
  rom[34739] = 16'hffff;
  rom[34740] = 16'hffff;
  rom[34741] = 16'hffff;
  rom[34742] = 16'hffff;
  rom[34743] = 16'hffff;
  rom[34744] = 16'hffff;
  rom[34745] = 16'hffff;
  rom[34746] = 16'hffff;
  rom[34747] = 16'hffff;
  rom[34748] = 16'hffff;
  rom[34749] = 16'hffff;
  rom[34750] = 16'hffff;
  rom[34751] = 16'hffff;
  rom[34752] = 16'hffff;
  rom[34753] = 16'hffff;
  rom[34754] = 16'hffff;
  rom[34755] = 16'hffff;
  rom[34756] = 16'hffff;
  rom[34757] = 16'hffff;
  rom[34758] = 16'hffff;
  rom[34759] = 16'hffff;
  rom[34760] = 16'hffff;
  rom[34761] = 16'hffff;
  rom[34762] = 16'hffff;
  rom[34763] = 16'hffff;
  rom[34764] = 16'hffff;
  rom[34765] = 16'hffff;
  rom[34766] = 16'hffff;
  rom[34767] = 16'hffff;
  rom[34768] = 16'hffff;
  rom[34769] = 16'hffff;
  rom[34770] = 16'hffff;
  rom[34771] = 16'hffff;
  rom[34772] = 16'hffff;
  rom[34773] = 16'hffff;
  rom[34774] = 16'hffff;
  rom[34775] = 16'hffff;
  rom[34776] = 16'hffff;
  rom[34777] = 16'hffff;
  rom[34778] = 16'hffff;
  rom[34779] = 16'hffff;
  rom[34780] = 16'hffff;
  rom[34781] = 16'hffff;
  rom[34782] = 16'hffff;
  rom[34783] = 16'hffff;
  rom[34784] = 16'hffff;
  rom[34785] = 16'hffff;
  rom[34786] = 16'hffff;
  rom[34787] = 16'hffff;
  rom[34788] = 16'hffff;
  rom[34789] = 16'hffff;
  rom[34790] = 16'hffff;
  rom[34791] = 16'hffff;
  rom[34792] = 16'hffff;
  rom[34793] = 16'hffff;
  rom[34794] = 16'hffff;
  rom[34795] = 16'hffff;
  rom[34796] = 16'hffff;
  rom[34797] = 16'hffff;
  rom[34798] = 16'hffff;
  rom[34799] = 16'hffff;
  rom[34800] = 16'hffff;
  rom[34801] = 16'hffff;
  rom[34802] = 16'hffff;
  rom[34803] = 16'hffff;
  rom[34804] = 16'hffff;
  rom[34805] = 16'hffff;
  rom[34806] = 16'hffff;
  rom[34807] = 16'hffff;
  rom[34808] = 16'hffff;
  rom[34809] = 16'hffff;
  rom[34810] = 16'hffff;
  rom[34811] = 16'hffff;
  rom[34812] = 16'hffff;
  rom[34813] = 16'hffff;
  rom[34814] = 16'hffff;
  rom[34815] = 16'hffff;
  rom[34816] = 16'hffff;
  rom[34817] = 16'hffff;
  rom[34818] = 16'hffff;
  rom[34819] = 16'hffff;
  rom[34820] = 16'hffff;
  rom[34821] = 16'hffff;
  rom[34822] = 16'hffff;
  rom[34823] = 16'hffff;
  rom[34824] = 16'hffff;
  rom[34825] = 16'hffff;
  rom[34826] = 16'hffff;
  rom[34827] = 16'hffff;
  rom[34828] = 16'hffff;
  rom[34829] = 16'hffff;
  rom[34830] = 16'hffff;
  rom[34831] = 16'hffff;
  rom[34832] = 16'hffff;
  rom[34833] = 16'hffff;
  rom[34834] = 16'hffff;
  rom[34835] = 16'hffff;
  rom[34836] = 16'hffff;
  rom[34837] = 16'hffff;
  rom[34838] = 16'hffff;
  rom[34839] = 16'hffff;
  rom[34840] = 16'hffff;
  rom[34841] = 16'hffff;
  rom[34842] = 16'hffff;
  rom[34843] = 16'hffff;
  rom[34844] = 16'hffff;
  rom[34845] = 16'hffff;
  rom[34846] = 16'hffff;
  rom[34847] = 16'hffff;
  rom[34848] = 16'hffff;
  rom[34849] = 16'hffff;
  rom[34850] = 16'hffff;
  rom[34851] = 16'hffff;
  rom[34852] = 16'hffff;
  rom[34853] = 16'hffff;
  rom[34854] = 16'hffff;
  rom[34855] = 16'hffff;
  rom[34856] = 16'hffff;
  rom[34857] = 16'hffff;
  rom[34858] = 16'hffff;
  rom[34859] = 16'hffff;
  rom[34860] = 16'hffff;
  rom[34861] = 16'hffff;
  rom[34862] = 16'hffff;
  rom[34863] = 16'hffff;
  rom[34864] = 16'hffff;
  rom[34865] = 16'hffff;
  rom[34866] = 16'hffff;
  rom[34867] = 16'hffff;
  rom[34868] = 16'hffff;
  rom[34869] = 16'hffff;
  rom[34870] = 16'hffff;
  rom[34871] = 16'hffff;
  rom[34872] = 16'hffdf;
  rom[34873] = 16'ha4ae;
  rom[34874] = 16'h7322;
  rom[34875] = 16'he68b;
  rom[34876] = 16'hf70a;
  rom[34877] = 16'hff0a;
  rom[34878] = 16'hff2a;
  rom[34879] = 16'hff28;
  rom[34880] = 16'hff08;
  rom[34881] = 16'hff28;
  rom[34882] = 16'hf708;
  rom[34883] = 16'hff28;
  rom[34884] = 16'hff08;
  rom[34885] = 16'hff28;
  rom[34886] = 16'hf708;
  rom[34887] = 16'hff28;
  rom[34888] = 16'hff08;
  rom[34889] = 16'hff28;
  rom[34890] = 16'hf728;
  rom[34891] = 16'hff29;
  rom[34892] = 16'hff09;
  rom[34893] = 16'hff28;
  rom[34894] = 16'hf708;
  rom[34895] = 16'hff0a;
  rom[34896] = 16'hf70a;
  rom[34897] = 16'hf72a;
  rom[34898] = 16'hde8a;
  rom[34899] = 16'h9403;
  rom[34900] = 16'hde8b;
  rom[34901] = 16'hef0b;
  rom[34902] = 16'hef09;
  rom[34903] = 16'hff49;
  rom[34904] = 16'hff09;
  rom[34905] = 16'hff2a;
  rom[34906] = 16'hf709;
  rom[34907] = 16'hff29;
  rom[34908] = 16'hff08;
  rom[34909] = 16'hff29;
  rom[34910] = 16'hff09;
  rom[34911] = 16'hff29;
  rom[34912] = 16'hff09;
  rom[34913] = 16'hff0b;
  rom[34914] = 16'hff2b;
  rom[34915] = 16'hf6e9;
  rom[34916] = 16'hf72c;
  rom[34917] = 16'hef0e;
  rom[34918] = 16'hd58b;
  rom[34919] = 16'h6961;
  rom[34920] = 16'hb245;
  rom[34921] = 16'hdaa8;
  rom[34922] = 16'hd288;
  rom[34923] = 16'hcaca;
  rom[34924] = 16'hfd54;
  rom[34925] = 16'hff5c;
  rom[34926] = 16'hfffe;
  rom[34927] = 16'hffff;
  rom[34928] = 16'hffff;
  rom[34929] = 16'hffff;
  rom[34930] = 16'hffff;
  rom[34931] = 16'hffff;
  rom[34932] = 16'hffff;
  rom[34933] = 16'hffff;
  rom[34934] = 16'hffff;
  rom[34935] = 16'hffff;
  rom[34936] = 16'hffff;
  rom[34937] = 16'hffff;
  rom[34938] = 16'hffff;
  rom[34939] = 16'hffff;
  rom[34940] = 16'hffff;
  rom[34941] = 16'hffff;
  rom[34942] = 16'hffff;
  rom[34943] = 16'hffff;
  rom[34944] = 16'hffff;
  rom[34945] = 16'hffff;
  rom[34946] = 16'hffff;
  rom[34947] = 16'hffff;
  rom[34948] = 16'hffff;
  rom[34949] = 16'hffff;
  rom[34950] = 16'hffff;
  rom[34951] = 16'hffff;
  rom[34952] = 16'hffff;
  rom[34953] = 16'hffff;
  rom[34954] = 16'hffff;
  rom[34955] = 16'hffff;
  rom[34956] = 16'hffff;
  rom[34957] = 16'hffff;
  rom[34958] = 16'hffff;
  rom[34959] = 16'hffff;
  rom[34960] = 16'hffff;
  rom[34961] = 16'hffff;
  rom[34962] = 16'hffff;
  rom[34963] = 16'hffff;
  rom[34964] = 16'hffff;
  rom[34965] = 16'hffff;
  rom[34966] = 16'hffff;
  rom[34967] = 16'hffff;
  rom[34968] = 16'hffff;
  rom[34969] = 16'hffff;
  rom[34970] = 16'hffff;
  rom[34971] = 16'hffff;
  rom[34972] = 16'hffff;
  rom[34973] = 16'hffff;
  rom[34974] = 16'hffff;
  rom[34975] = 16'hffff;
  rom[34976] = 16'hffff;
  rom[34977] = 16'hffff;
  rom[34978] = 16'hffff;
  rom[34979] = 16'hffff;
  rom[34980] = 16'hffff;
  rom[34981] = 16'hffff;
  rom[34982] = 16'hffff;
  rom[34983] = 16'hffff;
  rom[34984] = 16'hffff;
  rom[34985] = 16'hffff;
  rom[34986] = 16'hffff;
  rom[34987] = 16'hffff;
  rom[34988] = 16'hffff;
  rom[34989] = 16'hffff;
  rom[34990] = 16'hffff;
  rom[34991] = 16'hffff;
  rom[34992] = 16'hffff;
  rom[34993] = 16'hffff;
  rom[34994] = 16'hffff;
  rom[34995] = 16'hffff;
  rom[34996] = 16'hffff;
  rom[34997] = 16'hffff;
  rom[34998] = 16'hffff;
  rom[34999] = 16'hffff;
  rom[35000] = 16'hffff;
  rom[35001] = 16'hffff;
  rom[35002] = 16'hffff;
  rom[35003] = 16'hffff;
  rom[35004] = 16'hffff;
  rom[35005] = 16'hffff;
  rom[35006] = 16'hffff;
  rom[35007] = 16'hffff;
  rom[35008] = 16'hffff;
  rom[35009] = 16'hffff;
  rom[35010] = 16'hffff;
  rom[35011] = 16'hffff;
  rom[35012] = 16'hffff;
  rom[35013] = 16'hffff;
  rom[35014] = 16'hffff;
  rom[35015] = 16'hffff;
  rom[35016] = 16'hffff;
  rom[35017] = 16'hffff;
  rom[35018] = 16'hffff;
  rom[35019] = 16'hffff;
  rom[35020] = 16'hffff;
  rom[35021] = 16'hffff;
  rom[35022] = 16'hffff;
  rom[35023] = 16'hffff;
  rom[35024] = 16'hffff;
  rom[35025] = 16'hffff;
  rom[35026] = 16'hffff;
  rom[35027] = 16'hffff;
  rom[35028] = 16'hffff;
  rom[35029] = 16'hffff;
  rom[35030] = 16'hffff;
  rom[35031] = 16'hffff;
  rom[35032] = 16'hffff;
  rom[35033] = 16'hffff;
  rom[35034] = 16'hffff;
  rom[35035] = 16'hffff;
  rom[35036] = 16'hffff;
  rom[35037] = 16'hffff;
  rom[35038] = 16'hffff;
  rom[35039] = 16'hffff;
  rom[35040] = 16'hffff;
  rom[35041] = 16'hffff;
  rom[35042] = 16'hffff;
  rom[35043] = 16'hffff;
  rom[35044] = 16'hffff;
  rom[35045] = 16'hffff;
  rom[35046] = 16'hffff;
  rom[35047] = 16'hffff;
  rom[35048] = 16'hffff;
  rom[35049] = 16'hffff;
  rom[35050] = 16'hffff;
  rom[35051] = 16'hffff;
  rom[35052] = 16'hffff;
  rom[35053] = 16'hffff;
  rom[35054] = 16'hffff;
  rom[35055] = 16'hffff;
  rom[35056] = 16'hffff;
  rom[35057] = 16'hffff;
  rom[35058] = 16'hffff;
  rom[35059] = 16'hffff;
  rom[35060] = 16'hffff;
  rom[35061] = 16'hffff;
  rom[35062] = 16'hffff;
  rom[35063] = 16'hffff;
  rom[35064] = 16'hffff;
  rom[35065] = 16'hffff;
  rom[35066] = 16'hffff;
  rom[35067] = 16'hffff;
  rom[35068] = 16'hffff;
  rom[35069] = 16'hffff;
  rom[35070] = 16'hffff;
  rom[35071] = 16'hffff;
  rom[35072] = 16'hffff;
  rom[35073] = 16'hbdd3;
  rom[35074] = 16'h5261;
  rom[35075] = 16'hd62b;
  rom[35076] = 16'hff6c;
  rom[35077] = 16'hf709;
  rom[35078] = 16'hff4a;
  rom[35079] = 16'hf707;
  rom[35080] = 16'hff49;
  rom[35081] = 16'hff28;
  rom[35082] = 16'hff29;
  rom[35083] = 16'hff29;
  rom[35084] = 16'hff29;
  rom[35085] = 16'hff28;
  rom[35086] = 16'hff29;
  rom[35087] = 16'hff28;
  rom[35088] = 16'hff29;
  rom[35089] = 16'hff28;
  rom[35090] = 16'hf748;
  rom[35091] = 16'hf728;
  rom[35092] = 16'hff2a;
  rom[35093] = 16'hff28;
  rom[35094] = 16'hff29;
  rom[35095] = 16'hff0a;
  rom[35096] = 16'hff2b;
  rom[35097] = 16'hf72b;
  rom[35098] = 16'heeec;
  rom[35099] = 16'h9c84;
  rom[35100] = 16'hd649;
  rom[35101] = 16'hf72b;
  rom[35102] = 16'hf72b;
  rom[35103] = 16'hf70a;
  rom[35104] = 16'hff2a;
  rom[35105] = 16'hf709;
  rom[35106] = 16'hff2a;
  rom[35107] = 16'hf709;
  rom[35108] = 16'hff2a;
  rom[35109] = 16'hfee9;
  rom[35110] = 16'hff2b;
  rom[35111] = 16'hfeea;
  rom[35112] = 16'hff0b;
  rom[35113] = 16'hff0a;
  rom[35114] = 16'hf6ca;
  rom[35115] = 16'hff4c;
  rom[35116] = 16'hf6ce;
  rom[35117] = 16'hd56c;
  rom[35118] = 16'h8224;
  rom[35119] = 16'hbb08;
  rom[35120] = 16'hd2a8;
  rom[35121] = 16'hc268;
  rom[35122] = 16'hdbae;
  rom[35123] = 16'hf595;
  rom[35124] = 16'hff7e;
  rom[35125] = 16'hffbe;
  rom[35126] = 16'hffff;
  rom[35127] = 16'hffff;
  rom[35128] = 16'hffff;
  rom[35129] = 16'hffff;
  rom[35130] = 16'hffff;
  rom[35131] = 16'hffff;
  rom[35132] = 16'hffff;
  rom[35133] = 16'hffff;
  rom[35134] = 16'hffff;
  rom[35135] = 16'hffff;
  rom[35136] = 16'hffff;
  rom[35137] = 16'hffff;
  rom[35138] = 16'hffff;
  rom[35139] = 16'hffff;
  rom[35140] = 16'hffff;
  rom[35141] = 16'hffff;
  rom[35142] = 16'hffff;
  rom[35143] = 16'hffff;
  rom[35144] = 16'hffff;
  rom[35145] = 16'hffff;
  rom[35146] = 16'hffff;
  rom[35147] = 16'hffff;
  rom[35148] = 16'hffff;
  rom[35149] = 16'hffff;
  rom[35150] = 16'hffff;
  rom[35151] = 16'hffff;
  rom[35152] = 16'hffff;
  rom[35153] = 16'hffff;
  rom[35154] = 16'hffff;
  rom[35155] = 16'hffff;
  rom[35156] = 16'hffff;
  rom[35157] = 16'hffff;
  rom[35158] = 16'hffff;
  rom[35159] = 16'hffff;
  rom[35160] = 16'hffff;
  rom[35161] = 16'hffff;
  rom[35162] = 16'hffff;
  rom[35163] = 16'hffff;
  rom[35164] = 16'hffff;
  rom[35165] = 16'hffff;
  rom[35166] = 16'hffff;
  rom[35167] = 16'hffff;
  rom[35168] = 16'hffff;
  rom[35169] = 16'hffff;
  rom[35170] = 16'hffff;
  rom[35171] = 16'hffff;
  rom[35172] = 16'hffff;
  rom[35173] = 16'hffff;
  rom[35174] = 16'hffff;
  rom[35175] = 16'hffff;
  rom[35176] = 16'hffff;
  rom[35177] = 16'hffff;
  rom[35178] = 16'hffff;
  rom[35179] = 16'hffff;
  rom[35180] = 16'hffff;
  rom[35181] = 16'hffff;
  rom[35182] = 16'hffff;
  rom[35183] = 16'hffff;
  rom[35184] = 16'hffff;
  rom[35185] = 16'hffff;
  rom[35186] = 16'hffff;
  rom[35187] = 16'hffff;
  rom[35188] = 16'hffff;
  rom[35189] = 16'hffff;
  rom[35190] = 16'hffff;
  rom[35191] = 16'hffff;
  rom[35192] = 16'hffff;
  rom[35193] = 16'hffff;
  rom[35194] = 16'hffff;
  rom[35195] = 16'hffff;
  rom[35196] = 16'hffff;
  rom[35197] = 16'hffff;
  rom[35198] = 16'hffff;
  rom[35199] = 16'hffff;
  rom[35200] = 16'hffff;
  rom[35201] = 16'hffff;
  rom[35202] = 16'hffff;
  rom[35203] = 16'hffff;
  rom[35204] = 16'hffff;
  rom[35205] = 16'hffff;
  rom[35206] = 16'hffff;
  rom[35207] = 16'hffff;
  rom[35208] = 16'hffff;
  rom[35209] = 16'hffff;
  rom[35210] = 16'hffff;
  rom[35211] = 16'hffff;
  rom[35212] = 16'hffff;
  rom[35213] = 16'hffff;
  rom[35214] = 16'hffff;
  rom[35215] = 16'hffff;
  rom[35216] = 16'hffff;
  rom[35217] = 16'hffff;
  rom[35218] = 16'hffff;
  rom[35219] = 16'hffff;
  rom[35220] = 16'hffff;
  rom[35221] = 16'hffff;
  rom[35222] = 16'hffff;
  rom[35223] = 16'hffff;
  rom[35224] = 16'hffff;
  rom[35225] = 16'hffff;
  rom[35226] = 16'hffff;
  rom[35227] = 16'hffff;
  rom[35228] = 16'hffff;
  rom[35229] = 16'hffff;
  rom[35230] = 16'hffff;
  rom[35231] = 16'hffff;
  rom[35232] = 16'hffff;
  rom[35233] = 16'hffff;
  rom[35234] = 16'hffff;
  rom[35235] = 16'hffff;
  rom[35236] = 16'hffff;
  rom[35237] = 16'hffff;
  rom[35238] = 16'hffff;
  rom[35239] = 16'hffff;
  rom[35240] = 16'hffff;
  rom[35241] = 16'hffff;
  rom[35242] = 16'hffff;
  rom[35243] = 16'hffff;
  rom[35244] = 16'hffff;
  rom[35245] = 16'hffff;
  rom[35246] = 16'hffff;
  rom[35247] = 16'hffff;
  rom[35248] = 16'hffff;
  rom[35249] = 16'hffff;
  rom[35250] = 16'hffff;
  rom[35251] = 16'hffff;
  rom[35252] = 16'hffff;
  rom[35253] = 16'hffff;
  rom[35254] = 16'hffff;
  rom[35255] = 16'hffff;
  rom[35256] = 16'hffff;
  rom[35257] = 16'hffff;
  rom[35258] = 16'hffff;
  rom[35259] = 16'hffff;
  rom[35260] = 16'hffff;
  rom[35261] = 16'hffff;
  rom[35262] = 16'hffff;
  rom[35263] = 16'hffff;
  rom[35264] = 16'hffff;
  rom[35265] = 16'hffff;
  rom[35266] = 16'hffff;
  rom[35267] = 16'hffff;
  rom[35268] = 16'hffff;
  rom[35269] = 16'hffff;
  rom[35270] = 16'hffdf;
  rom[35271] = 16'hffff;
  rom[35272] = 16'hfffe;
  rom[35273] = 16'hded8;
  rom[35274] = 16'h5283;
  rom[35275] = 16'hce2c;
  rom[35276] = 16'hf74b;
  rom[35277] = 16'heee9;
  rom[35278] = 16'hf708;
  rom[35279] = 16'hf708;
  rom[35280] = 16'hf728;
  rom[35281] = 16'hff28;
  rom[35282] = 16'hff08;
  rom[35283] = 16'hff49;
  rom[35284] = 16'hf708;
  rom[35285] = 16'hff28;
  rom[35286] = 16'hff08;
  rom[35287] = 16'hff28;
  rom[35288] = 16'hf708;
  rom[35289] = 16'hff28;
  rom[35290] = 16'hf727;
  rom[35291] = 16'hf748;
  rom[35292] = 16'hf708;
  rom[35293] = 16'hff29;
  rom[35294] = 16'hff09;
  rom[35295] = 16'hff2a;
  rom[35296] = 16'hf72a;
  rom[35297] = 16'hef0a;
  rom[35298] = 16'he6cb;
  rom[35299] = 16'h9ca5;
  rom[35300] = 16'had04;
  rom[35301] = 16'hf72c;
  rom[35302] = 16'heee9;
  rom[35303] = 16'hff2a;
  rom[35304] = 16'hf749;
  rom[35305] = 16'hff29;
  rom[35306] = 16'hf708;
  rom[35307] = 16'hff49;
  rom[35308] = 16'hff08;
  rom[35309] = 16'hff09;
  rom[35310] = 16'hff0a;
  rom[35311] = 16'hff2b;
  rom[35312] = 16'hff0b;
  rom[35313] = 16'hf72b;
  rom[35314] = 16'hf70c;
  rom[35315] = 16'hf6ce;
  rom[35316] = 16'hbca9;
  rom[35317] = 16'h6942;
  rom[35318] = 16'hb2a8;
  rom[35319] = 16'hb248;
  rom[35320] = 16'hbaaa;
  rom[35321] = 16'hecb2;
  rom[35322] = 16'hfe59;
  rom[35323] = 16'hff9e;
  rom[35324] = 16'hffbe;
  rom[35325] = 16'hffff;
  rom[35326] = 16'hffff;
  rom[35327] = 16'hffff;
  rom[35328] = 16'hffdf;
  rom[35329] = 16'hffff;
  rom[35330] = 16'hffff;
  rom[35331] = 16'hffff;
  rom[35332] = 16'hffff;
  rom[35333] = 16'hffff;
  rom[35334] = 16'hffff;
  rom[35335] = 16'hffff;
  rom[35336] = 16'hffff;
  rom[35337] = 16'hffff;
  rom[35338] = 16'hffff;
  rom[35339] = 16'hffff;
  rom[35340] = 16'hffff;
  rom[35341] = 16'hffff;
  rom[35342] = 16'hffff;
  rom[35343] = 16'hffff;
  rom[35344] = 16'hffff;
  rom[35345] = 16'hffff;
  rom[35346] = 16'hffff;
  rom[35347] = 16'hffff;
  rom[35348] = 16'hffff;
  rom[35349] = 16'hffff;
  rom[35350] = 16'hffff;
  rom[35351] = 16'hffff;
  rom[35352] = 16'hffff;
  rom[35353] = 16'hffff;
  rom[35354] = 16'hffff;
  rom[35355] = 16'hffff;
  rom[35356] = 16'hffff;
  rom[35357] = 16'hffff;
  rom[35358] = 16'hffff;
  rom[35359] = 16'hffff;
  rom[35360] = 16'hffff;
  rom[35361] = 16'hffff;
  rom[35362] = 16'hffff;
  rom[35363] = 16'hffff;
  rom[35364] = 16'hffff;
  rom[35365] = 16'hffff;
  rom[35366] = 16'hffff;
  rom[35367] = 16'hffff;
  rom[35368] = 16'hffff;
  rom[35369] = 16'hffff;
  rom[35370] = 16'hffff;
  rom[35371] = 16'hffff;
  rom[35372] = 16'hffff;
  rom[35373] = 16'hffff;
  rom[35374] = 16'hffff;
  rom[35375] = 16'hffff;
  rom[35376] = 16'hffff;
  rom[35377] = 16'hffff;
  rom[35378] = 16'hffff;
  rom[35379] = 16'hffff;
  rom[35380] = 16'hffff;
  rom[35381] = 16'hffff;
  rom[35382] = 16'hffff;
  rom[35383] = 16'hffff;
  rom[35384] = 16'hffff;
  rom[35385] = 16'hffff;
  rom[35386] = 16'hffff;
  rom[35387] = 16'hffff;
  rom[35388] = 16'hffff;
  rom[35389] = 16'hffff;
  rom[35390] = 16'hffff;
  rom[35391] = 16'hffff;
  rom[35392] = 16'hffff;
  rom[35393] = 16'hffff;
  rom[35394] = 16'hffff;
  rom[35395] = 16'hffff;
  rom[35396] = 16'hffff;
  rom[35397] = 16'hffff;
  rom[35398] = 16'hffff;
  rom[35399] = 16'hffff;
  rom[35400] = 16'hffff;
  rom[35401] = 16'hffff;
  rom[35402] = 16'hffff;
  rom[35403] = 16'hffff;
  rom[35404] = 16'hffff;
  rom[35405] = 16'hffff;
  rom[35406] = 16'hffff;
  rom[35407] = 16'hffff;
  rom[35408] = 16'hffff;
  rom[35409] = 16'hffff;
  rom[35410] = 16'hffff;
  rom[35411] = 16'hffff;
  rom[35412] = 16'hffff;
  rom[35413] = 16'hffff;
  rom[35414] = 16'hffff;
  rom[35415] = 16'hffff;
  rom[35416] = 16'hffff;
  rom[35417] = 16'hffff;
  rom[35418] = 16'hffff;
  rom[35419] = 16'hffff;
  rom[35420] = 16'hffff;
  rom[35421] = 16'hffff;
  rom[35422] = 16'hffff;
  rom[35423] = 16'hffff;
  rom[35424] = 16'hffff;
  rom[35425] = 16'hffff;
  rom[35426] = 16'hffff;
  rom[35427] = 16'hffff;
  rom[35428] = 16'hffff;
  rom[35429] = 16'hffff;
  rom[35430] = 16'hffff;
  rom[35431] = 16'hffff;
  rom[35432] = 16'hffff;
  rom[35433] = 16'hffff;
  rom[35434] = 16'hffff;
  rom[35435] = 16'hffff;
  rom[35436] = 16'hffff;
  rom[35437] = 16'hffff;
  rom[35438] = 16'hffff;
  rom[35439] = 16'hffff;
  rom[35440] = 16'hffff;
  rom[35441] = 16'hffff;
  rom[35442] = 16'hffff;
  rom[35443] = 16'hffff;
  rom[35444] = 16'hffff;
  rom[35445] = 16'hffff;
  rom[35446] = 16'hffff;
  rom[35447] = 16'hffff;
  rom[35448] = 16'hffff;
  rom[35449] = 16'hffff;
  rom[35450] = 16'hffff;
  rom[35451] = 16'hffff;
  rom[35452] = 16'hffff;
  rom[35453] = 16'hffff;
  rom[35454] = 16'hffff;
  rom[35455] = 16'hffff;
  rom[35456] = 16'hffff;
  rom[35457] = 16'hffff;
  rom[35458] = 16'hffff;
  rom[35459] = 16'hffff;
  rom[35460] = 16'hffff;
  rom[35461] = 16'hffff;
  rom[35462] = 16'hffff;
  rom[35463] = 16'hffff;
  rom[35464] = 16'hffff;
  rom[35465] = 16'hffff;
  rom[35466] = 16'hffff;
  rom[35467] = 16'hffff;
  rom[35468] = 16'hffff;
  rom[35469] = 16'hffff;
  rom[35470] = 16'hffff;
  rom[35471] = 16'hffff;
  rom[35472] = 16'hffff;
  rom[35473] = 16'hfffe;
  rom[35474] = 16'h7328;
  rom[35475] = 16'h94a7;
  rom[35476] = 16'hef4d;
  rom[35477] = 16'hf72a;
  rom[35478] = 16'hf729;
  rom[35479] = 16'hff28;
  rom[35480] = 16'hff29;
  rom[35481] = 16'hff28;
  rom[35482] = 16'hff29;
  rom[35483] = 16'hff29;
  rom[35484] = 16'hff29;
  rom[35485] = 16'hff28;
  rom[35486] = 16'hff29;
  rom[35487] = 16'hff28;
  rom[35488] = 16'hff29;
  rom[35489] = 16'hff28;
  rom[35490] = 16'hff48;
  rom[35491] = 16'hf727;
  rom[35492] = 16'hff29;
  rom[35493] = 16'hff09;
  rom[35494] = 16'hff0a;
  rom[35495] = 16'hff29;
  rom[35496] = 16'hf729;
  rom[35497] = 16'hf72a;
  rom[35498] = 16'hff6d;
  rom[35499] = 16'hbda8;
  rom[35500] = 16'h7340;
  rom[35501] = 16'hde6a;
  rom[35502] = 16'hf70c;
  rom[35503] = 16'hf6ea;
  rom[35504] = 16'hff2a;
  rom[35505] = 16'hff49;
  rom[35506] = 16'hff29;
  rom[35507] = 16'hff28;
  rom[35508] = 16'hff29;
  rom[35509] = 16'hff29;
  rom[35510] = 16'hf70a;
  rom[35511] = 16'hff2b;
  rom[35512] = 16'hf70b;
  rom[35513] = 16'hf70c;
  rom[35514] = 16'heead;
  rom[35515] = 16'ha427;
  rom[35516] = 16'h7a64;
  rom[35517] = 16'ha2c8;
  rom[35518] = 16'hc34c;
  rom[35519] = 16'hd3ef;
  rom[35520] = 16'hf5b6;
  rom[35521] = 16'hff3c;
  rom[35522] = 16'hffdf;
  rom[35523] = 16'hffdf;
  rom[35524] = 16'hffff;
  rom[35525] = 16'hffff;
  rom[35526] = 16'hffff;
  rom[35527] = 16'hffff;
  rom[35528] = 16'hffff;
  rom[35529] = 16'hffff;
  rom[35530] = 16'hffff;
  rom[35531] = 16'hffff;
  rom[35532] = 16'hffff;
  rom[35533] = 16'hffff;
  rom[35534] = 16'hffff;
  rom[35535] = 16'hffff;
  rom[35536] = 16'hffff;
  rom[35537] = 16'hffff;
  rom[35538] = 16'hffff;
  rom[35539] = 16'hffff;
  rom[35540] = 16'hffff;
  rom[35541] = 16'hffff;
  rom[35542] = 16'hffff;
  rom[35543] = 16'hffff;
  rom[35544] = 16'hffff;
  rom[35545] = 16'hffff;
  rom[35546] = 16'hffff;
  rom[35547] = 16'hffff;
  rom[35548] = 16'hffff;
  rom[35549] = 16'hffff;
  rom[35550] = 16'hffff;
  rom[35551] = 16'hffff;
  rom[35552] = 16'hffff;
  rom[35553] = 16'hffff;
  rom[35554] = 16'hffff;
  rom[35555] = 16'hffff;
  rom[35556] = 16'hffff;
  rom[35557] = 16'hffff;
  rom[35558] = 16'hffff;
  rom[35559] = 16'hffff;
  rom[35560] = 16'hffff;
  rom[35561] = 16'hffff;
  rom[35562] = 16'hffff;
  rom[35563] = 16'hffff;
  rom[35564] = 16'hffff;
  rom[35565] = 16'hffff;
  rom[35566] = 16'hffff;
  rom[35567] = 16'hffff;
  rom[35568] = 16'hffff;
  rom[35569] = 16'hffff;
  rom[35570] = 16'hffff;
  rom[35571] = 16'hffff;
  rom[35572] = 16'hffff;
  rom[35573] = 16'hffff;
  rom[35574] = 16'hffff;
  rom[35575] = 16'hffff;
  rom[35576] = 16'hffff;
  rom[35577] = 16'hffff;
  rom[35578] = 16'hffff;
  rom[35579] = 16'hffff;
  rom[35580] = 16'hffff;
  rom[35581] = 16'hffff;
  rom[35582] = 16'hffff;
  rom[35583] = 16'hffff;
  rom[35584] = 16'hffff;
  rom[35585] = 16'hffff;
  rom[35586] = 16'hffff;
  rom[35587] = 16'hffff;
  rom[35588] = 16'hffff;
  rom[35589] = 16'hffff;
  rom[35590] = 16'hffff;
  rom[35591] = 16'hffff;
  rom[35592] = 16'hffff;
  rom[35593] = 16'hffff;
  rom[35594] = 16'hffff;
  rom[35595] = 16'hffff;
  rom[35596] = 16'hffff;
  rom[35597] = 16'hffff;
  rom[35598] = 16'hffff;
  rom[35599] = 16'hffff;
  rom[35600] = 16'hffff;
  rom[35601] = 16'hffff;
  rom[35602] = 16'hffff;
  rom[35603] = 16'hffff;
  rom[35604] = 16'hffff;
  rom[35605] = 16'hffff;
  rom[35606] = 16'hffff;
  rom[35607] = 16'hffff;
  rom[35608] = 16'hffff;
  rom[35609] = 16'hffff;
  rom[35610] = 16'hffff;
  rom[35611] = 16'hffff;
  rom[35612] = 16'hffff;
  rom[35613] = 16'hffff;
  rom[35614] = 16'hffff;
  rom[35615] = 16'hffff;
  rom[35616] = 16'hffff;
  rom[35617] = 16'hffff;
  rom[35618] = 16'hffff;
  rom[35619] = 16'hffff;
  rom[35620] = 16'hffff;
  rom[35621] = 16'hffff;
  rom[35622] = 16'hffff;
  rom[35623] = 16'hffff;
  rom[35624] = 16'hffff;
  rom[35625] = 16'hffff;
  rom[35626] = 16'hffff;
  rom[35627] = 16'hffff;
  rom[35628] = 16'hffff;
  rom[35629] = 16'hffff;
  rom[35630] = 16'hffff;
  rom[35631] = 16'hffff;
  rom[35632] = 16'hffff;
  rom[35633] = 16'hffff;
  rom[35634] = 16'hffff;
  rom[35635] = 16'hffff;
  rom[35636] = 16'hffff;
  rom[35637] = 16'hffff;
  rom[35638] = 16'hffff;
  rom[35639] = 16'hffff;
  rom[35640] = 16'hffff;
  rom[35641] = 16'hffff;
  rom[35642] = 16'hffff;
  rom[35643] = 16'hffff;
  rom[35644] = 16'hffff;
  rom[35645] = 16'hffff;
  rom[35646] = 16'hffff;
  rom[35647] = 16'hffff;
  rom[35648] = 16'hffff;
  rom[35649] = 16'hffff;
  rom[35650] = 16'hffff;
  rom[35651] = 16'hffff;
  rom[35652] = 16'hffff;
  rom[35653] = 16'hffff;
  rom[35654] = 16'hffff;
  rom[35655] = 16'hffff;
  rom[35656] = 16'hffff;
  rom[35657] = 16'hffff;
  rom[35658] = 16'hffff;
  rom[35659] = 16'hffff;
  rom[35660] = 16'hffff;
  rom[35661] = 16'hffff;
  rom[35662] = 16'hffff;
  rom[35663] = 16'hffff;
  rom[35664] = 16'hffff;
  rom[35665] = 16'hffff;
  rom[35666] = 16'hffff;
  rom[35667] = 16'hffff;
  rom[35668] = 16'hffff;
  rom[35669] = 16'hffff;
  rom[35670] = 16'hffff;
  rom[35671] = 16'hffff;
  rom[35672] = 16'hffdf;
  rom[35673] = 16'hffff;
  rom[35674] = 16'h9c6e;
  rom[35675] = 16'h83c6;
  rom[35676] = 16'hef2d;
  rom[35677] = 16'hff6b;
  rom[35678] = 16'heee8;
  rom[35679] = 16'hff49;
  rom[35680] = 16'hff08;
  rom[35681] = 16'hff28;
  rom[35682] = 16'hf708;
  rom[35683] = 16'hf729;
  rom[35684] = 16'hff29;
  rom[35685] = 16'hff29;
  rom[35686] = 16'hf709;
  rom[35687] = 16'hff29;
  rom[35688] = 16'hff08;
  rom[35689] = 16'hff28;
  rom[35690] = 16'hf728;
  rom[35691] = 16'hf748;
  rom[35692] = 16'hff09;
  rom[35693] = 16'hff0a;
  rom[35694] = 16'hf709;
  rom[35695] = 16'hff28;
  rom[35696] = 16'hf728;
  rom[35697] = 16'hff4a;
  rom[35698] = 16'heeca;
  rom[35699] = 16'he6ac;
  rom[35700] = 16'h83a3;
  rom[35701] = 16'hac85;
  rom[35702] = 16'hf6ac;
  rom[35703] = 16'hf70c;
  rom[35704] = 16'hff0b;
  rom[35705] = 16'hff2a;
  rom[35706] = 16'hf749;
  rom[35707] = 16'hff4a;
  rom[35708] = 16'hf72a;
  rom[35709] = 16'hf70a;
  rom[35710] = 16'hf70b;
  rom[35711] = 16'hf72d;
  rom[35712] = 16'heeed;
  rom[35713] = 16'hcd8a;
  rom[35714] = 16'h7b23;
  rom[35715] = 16'h7ac5;
  rom[35716] = 16'h9b8b;
  rom[35717] = 16'hcc91;
  rom[35718] = 16'hee17;
  rom[35719] = 16'hfeba;
  rom[35720] = 16'hff9d;
  rom[35721] = 16'hffff;
  rom[35722] = 16'hffdf;
  rom[35723] = 16'hffff;
  rom[35724] = 16'hffff;
  rom[35725] = 16'hffff;
  rom[35726] = 16'hffdf;
  rom[35727] = 16'hffff;
  rom[35728] = 16'hffff;
  rom[35729] = 16'hffff;
  rom[35730] = 16'hffff;
  rom[35731] = 16'hffff;
  rom[35732] = 16'hffff;
  rom[35733] = 16'hffff;
  rom[35734] = 16'hffff;
  rom[35735] = 16'hffff;
  rom[35736] = 16'hffff;
  rom[35737] = 16'hffff;
  rom[35738] = 16'hffff;
  rom[35739] = 16'hffff;
  rom[35740] = 16'hffff;
  rom[35741] = 16'hffff;
  rom[35742] = 16'hffff;
  rom[35743] = 16'hffff;
  rom[35744] = 16'hffff;
  rom[35745] = 16'hffff;
  rom[35746] = 16'hffff;
  rom[35747] = 16'hffff;
  rom[35748] = 16'hffff;
  rom[35749] = 16'hffff;
  rom[35750] = 16'hffff;
  rom[35751] = 16'hffff;
  rom[35752] = 16'hffff;
  rom[35753] = 16'hffff;
  rom[35754] = 16'hffff;
  rom[35755] = 16'hffff;
  rom[35756] = 16'hffff;
  rom[35757] = 16'hffff;
  rom[35758] = 16'hffff;
  rom[35759] = 16'hffff;
  rom[35760] = 16'hffff;
  rom[35761] = 16'hffff;
  rom[35762] = 16'hffff;
  rom[35763] = 16'hffff;
  rom[35764] = 16'hffff;
  rom[35765] = 16'hffff;
  rom[35766] = 16'hffff;
  rom[35767] = 16'hffff;
  rom[35768] = 16'hffff;
  rom[35769] = 16'hffff;
  rom[35770] = 16'hffff;
  rom[35771] = 16'hffff;
  rom[35772] = 16'hffff;
  rom[35773] = 16'hffff;
  rom[35774] = 16'hffff;
  rom[35775] = 16'hffff;
  rom[35776] = 16'hffff;
  rom[35777] = 16'hffff;
  rom[35778] = 16'hffff;
  rom[35779] = 16'hffff;
  rom[35780] = 16'hffff;
  rom[35781] = 16'hffff;
  rom[35782] = 16'hffff;
  rom[35783] = 16'hffff;
  rom[35784] = 16'hffff;
  rom[35785] = 16'hffff;
  rom[35786] = 16'hffff;
  rom[35787] = 16'hffff;
  rom[35788] = 16'hffff;
  rom[35789] = 16'hffff;
  rom[35790] = 16'hffff;
  rom[35791] = 16'hffff;
  rom[35792] = 16'hffff;
  rom[35793] = 16'hffff;
  rom[35794] = 16'hffff;
  rom[35795] = 16'hffff;
  rom[35796] = 16'hffff;
  rom[35797] = 16'hffff;
  rom[35798] = 16'hffff;
  rom[35799] = 16'hffff;
  rom[35800] = 16'hffff;
  rom[35801] = 16'hffff;
  rom[35802] = 16'hffff;
  rom[35803] = 16'hffff;
  rom[35804] = 16'hffff;
  rom[35805] = 16'hffff;
  rom[35806] = 16'hffff;
  rom[35807] = 16'hffff;
  rom[35808] = 16'hffff;
  rom[35809] = 16'hffff;
  rom[35810] = 16'hffff;
  rom[35811] = 16'hffff;
  rom[35812] = 16'hffff;
  rom[35813] = 16'hffff;
  rom[35814] = 16'hffff;
  rom[35815] = 16'hffff;
  rom[35816] = 16'hffff;
  rom[35817] = 16'hffff;
  rom[35818] = 16'hffff;
  rom[35819] = 16'hffff;
  rom[35820] = 16'hffff;
  rom[35821] = 16'hffff;
  rom[35822] = 16'hffff;
  rom[35823] = 16'hffff;
  rom[35824] = 16'hffff;
  rom[35825] = 16'hffff;
  rom[35826] = 16'hffff;
  rom[35827] = 16'hffff;
  rom[35828] = 16'hffff;
  rom[35829] = 16'hffff;
  rom[35830] = 16'hffff;
  rom[35831] = 16'hffff;
  rom[35832] = 16'hffff;
  rom[35833] = 16'hffff;
  rom[35834] = 16'hffff;
  rom[35835] = 16'hffff;
  rom[35836] = 16'hffff;
  rom[35837] = 16'hffff;
  rom[35838] = 16'hffff;
  rom[35839] = 16'hffff;
  rom[35840] = 16'hffff;
  rom[35841] = 16'hffff;
  rom[35842] = 16'hffff;
  rom[35843] = 16'hffff;
  rom[35844] = 16'hffff;
  rom[35845] = 16'hffff;
  rom[35846] = 16'hffff;
  rom[35847] = 16'hffff;
  rom[35848] = 16'hffff;
  rom[35849] = 16'hffff;
  rom[35850] = 16'hffff;
  rom[35851] = 16'hffff;
  rom[35852] = 16'hffff;
  rom[35853] = 16'hffff;
  rom[35854] = 16'hffff;
  rom[35855] = 16'hffff;
  rom[35856] = 16'hffff;
  rom[35857] = 16'hffff;
  rom[35858] = 16'hffff;
  rom[35859] = 16'hffff;
  rom[35860] = 16'hffff;
  rom[35861] = 16'hffff;
  rom[35862] = 16'hffff;
  rom[35863] = 16'hffff;
  rom[35864] = 16'hffff;
  rom[35865] = 16'hffff;
  rom[35866] = 16'hffff;
  rom[35867] = 16'hffff;
  rom[35868] = 16'hffff;
  rom[35869] = 16'hffff;
  rom[35870] = 16'hffff;
  rom[35871] = 16'hffff;
  rom[35872] = 16'hffff;
  rom[35873] = 16'hffff;
  rom[35874] = 16'hde98;
  rom[35875] = 16'h7325;
  rom[35876] = 16'he6ad;
  rom[35877] = 16'heee9;
  rom[35878] = 16'hff69;
  rom[35879] = 16'hff49;
  rom[35880] = 16'hff29;
  rom[35881] = 16'hff29;
  rom[35882] = 16'hff29;
  rom[35883] = 16'hf708;
  rom[35884] = 16'hff4a;
  rom[35885] = 16'hff29;
  rom[35886] = 16'hff29;
  rom[35887] = 16'hff28;
  rom[35888] = 16'hff29;
  rom[35889] = 16'hff28;
  rom[35890] = 16'hff49;
  rom[35891] = 16'hff28;
  rom[35892] = 16'hff0a;
  rom[35893] = 16'hff0b;
  rom[35894] = 16'hff2a;
  rom[35895] = 16'hff27;
  rom[35896] = 16'hff48;
  rom[35897] = 16'hff29;
  rom[35898] = 16'hf72c;
  rom[35899] = 16'hf70d;
  rom[35900] = 16'hbd2a;
  rom[35901] = 16'h6200;
  rom[35902] = 16'hbcc8;
  rom[35903] = 16'hee8d;
  rom[35904] = 16'hfecd;
  rom[35905] = 16'hf6cc;
  rom[35906] = 16'hf70c;
  rom[35907] = 16'hef0b;
  rom[35908] = 16'hff4d;
  rom[35909] = 16'hef0d;
  rom[35910] = 16'he6cd;
  rom[35911] = 16'hc60b;
  rom[35912] = 16'h9467;
  rom[35913] = 16'h6ae3;
  rom[35914] = 16'h93ea;
  rom[35915] = 16'hcd73;
  rom[35916] = 16'hfeba;
  rom[35917] = 16'hff3c;
  rom[35918] = 16'hffbd;
  rom[35919] = 16'hfffe;
  rom[35920] = 16'hfffe;
  rom[35921] = 16'hffff;
  rom[35922] = 16'hffff;
  rom[35923] = 16'hffdf;
  rom[35924] = 16'hffff;
  rom[35925] = 16'hffff;
  rom[35926] = 16'hffff;
  rom[35927] = 16'hffff;
  rom[35928] = 16'hffff;
  rom[35929] = 16'hffff;
  rom[35930] = 16'hffff;
  rom[35931] = 16'hffff;
  rom[35932] = 16'hffff;
  rom[35933] = 16'hffff;
  rom[35934] = 16'hffff;
  rom[35935] = 16'hffff;
  rom[35936] = 16'hffff;
  rom[35937] = 16'hffff;
  rom[35938] = 16'hffff;
  rom[35939] = 16'hffff;
  rom[35940] = 16'hffff;
  rom[35941] = 16'hffff;
  rom[35942] = 16'hffff;
  rom[35943] = 16'hffff;
  rom[35944] = 16'hffff;
  rom[35945] = 16'hffff;
  rom[35946] = 16'hffff;
  rom[35947] = 16'hffff;
  rom[35948] = 16'hffff;
  rom[35949] = 16'hffff;
  rom[35950] = 16'hffff;
  rom[35951] = 16'hffff;
  rom[35952] = 16'hffff;
  rom[35953] = 16'hffff;
  rom[35954] = 16'hffff;
  rom[35955] = 16'hffff;
  rom[35956] = 16'hffff;
  rom[35957] = 16'hffff;
  rom[35958] = 16'hffff;
  rom[35959] = 16'hffff;
  rom[35960] = 16'hffff;
  rom[35961] = 16'hffff;
  rom[35962] = 16'hffff;
  rom[35963] = 16'hffff;
  rom[35964] = 16'hffff;
  rom[35965] = 16'hffff;
  rom[35966] = 16'hffff;
  rom[35967] = 16'hffff;
  rom[35968] = 16'hffff;
  rom[35969] = 16'hffff;
  rom[35970] = 16'hffff;
  rom[35971] = 16'hffff;
  rom[35972] = 16'hffff;
  rom[35973] = 16'hffff;
  rom[35974] = 16'hffff;
  rom[35975] = 16'hffff;
  rom[35976] = 16'hffff;
  rom[35977] = 16'hffff;
  rom[35978] = 16'hffff;
  rom[35979] = 16'hffff;
  rom[35980] = 16'hffff;
  rom[35981] = 16'hffff;
  rom[35982] = 16'hffff;
  rom[35983] = 16'hffff;
  rom[35984] = 16'hffff;
  rom[35985] = 16'hffff;
  rom[35986] = 16'hffff;
  rom[35987] = 16'hffff;
  rom[35988] = 16'hffff;
  rom[35989] = 16'hffff;
  rom[35990] = 16'hffff;
  rom[35991] = 16'hffff;
  rom[35992] = 16'hffff;
  rom[35993] = 16'hffff;
  rom[35994] = 16'hffff;
  rom[35995] = 16'hffff;
  rom[35996] = 16'hffff;
  rom[35997] = 16'hffff;
  rom[35998] = 16'hffff;
  rom[35999] = 16'hffff;
  rom[36000] = 16'hffff;
  rom[36001] = 16'hffff;
  rom[36002] = 16'hffff;
  rom[36003] = 16'hffff;
  rom[36004] = 16'hffff;
  rom[36005] = 16'hffff;
  rom[36006] = 16'hffff;
  rom[36007] = 16'hffff;
  rom[36008] = 16'hffff;
  rom[36009] = 16'hffff;
  rom[36010] = 16'hffff;
  rom[36011] = 16'hffff;
  rom[36012] = 16'hffff;
  rom[36013] = 16'hffff;
  rom[36014] = 16'hffff;
  rom[36015] = 16'hffff;
  rom[36016] = 16'hffff;
  rom[36017] = 16'hffff;
  rom[36018] = 16'hffff;
  rom[36019] = 16'hffff;
  rom[36020] = 16'hffff;
  rom[36021] = 16'hffff;
  rom[36022] = 16'hffff;
  rom[36023] = 16'hffff;
  rom[36024] = 16'hffff;
  rom[36025] = 16'hffff;
  rom[36026] = 16'hffff;
  rom[36027] = 16'hffff;
  rom[36028] = 16'hffff;
  rom[36029] = 16'hffff;
  rom[36030] = 16'hffff;
  rom[36031] = 16'hffff;
  rom[36032] = 16'hffff;
  rom[36033] = 16'hffff;
  rom[36034] = 16'hffff;
  rom[36035] = 16'hffff;
  rom[36036] = 16'hffff;
  rom[36037] = 16'hffff;
  rom[36038] = 16'hffff;
  rom[36039] = 16'hffff;
  rom[36040] = 16'hffff;
  rom[36041] = 16'hffff;
  rom[36042] = 16'hffff;
  rom[36043] = 16'hffff;
  rom[36044] = 16'hffff;
  rom[36045] = 16'hffff;
  rom[36046] = 16'hffff;
  rom[36047] = 16'hffff;
  rom[36048] = 16'hffff;
  rom[36049] = 16'hffff;
  rom[36050] = 16'hffff;
  rom[36051] = 16'hffff;
  rom[36052] = 16'hffff;
  rom[36053] = 16'hffff;
  rom[36054] = 16'hffff;
  rom[36055] = 16'hffff;
  rom[36056] = 16'hffff;
  rom[36057] = 16'hffff;
  rom[36058] = 16'hffff;
  rom[36059] = 16'hffff;
  rom[36060] = 16'hffff;
  rom[36061] = 16'hffff;
  rom[36062] = 16'hffff;
  rom[36063] = 16'hffff;
  rom[36064] = 16'hffff;
  rom[36065] = 16'hffff;
  rom[36066] = 16'hffff;
  rom[36067] = 16'hffff;
  rom[36068] = 16'hffff;
  rom[36069] = 16'hffff;
  rom[36070] = 16'hffff;
  rom[36071] = 16'hffff;
  rom[36072] = 16'hffff;
  rom[36073] = 16'hffff;
  rom[36074] = 16'hf77c;
  rom[36075] = 16'h6b05;
  rom[36076] = 16'hcdea;
  rom[36077] = 16'hf72b;
  rom[36078] = 16'hf708;
  rom[36079] = 16'hff29;
  rom[36080] = 16'hff09;
  rom[36081] = 16'hf709;
  rom[36082] = 16'hff29;
  rom[36083] = 16'hff28;
  rom[36084] = 16'hf728;
  rom[36085] = 16'hff28;
  rom[36086] = 16'hff08;
  rom[36087] = 16'hff28;
  rom[36088] = 16'hf708;
  rom[36089] = 16'hff29;
  rom[36090] = 16'hff08;
  rom[36091] = 16'hff29;
  rom[36092] = 16'hf709;
  rom[36093] = 16'hff0a;
  rom[36094] = 16'hff09;
  rom[36095] = 16'hff27;
  rom[36096] = 16'hf727;
  rom[36097] = 16'hff08;
  rom[36098] = 16'hf709;
  rom[36099] = 16'hff2d;
  rom[36100] = 16'ha447;
  rom[36101] = 16'h6201;
  rom[36102] = 16'h6a41;
  rom[36103] = 16'h9385;
  rom[36104] = 16'hb4c9;
  rom[36105] = 16'hd5ed;
  rom[36106] = 16'hd60d;
  rom[36107] = 16'hcded;
  rom[36108] = 16'hbd8b;
  rom[36109] = 16'ha50a;
  rom[36110] = 16'h8407;
  rom[36111] = 16'h8408;
  rom[36112] = 16'ha50e;
  rom[36113] = 16'he6b7;
  rom[36114] = 16'heefa;
  rom[36115] = 16'hff7d;
  rom[36116] = 16'hff9e;
  rom[36117] = 16'hffde;
  rom[36118] = 16'hffde;
  rom[36119] = 16'hf7de;
  rom[36120] = 16'hf7fe;
  rom[36121] = 16'hffff;
  rom[36122] = 16'hffff;
  rom[36123] = 16'hffff;
  rom[36124] = 16'hffde;
  rom[36125] = 16'hffff;
  rom[36126] = 16'hffff;
  rom[36127] = 16'hffff;
  rom[36128] = 16'hffff;
  rom[36129] = 16'hffff;
  rom[36130] = 16'hffff;
  rom[36131] = 16'hffff;
  rom[36132] = 16'hffff;
  rom[36133] = 16'hffff;
  rom[36134] = 16'hffff;
  rom[36135] = 16'hffff;
  rom[36136] = 16'hffff;
  rom[36137] = 16'hffff;
  rom[36138] = 16'hffff;
  rom[36139] = 16'hffff;
  rom[36140] = 16'hffff;
  rom[36141] = 16'hffff;
  rom[36142] = 16'hffff;
  rom[36143] = 16'hffff;
  rom[36144] = 16'hffff;
  rom[36145] = 16'hffff;
  rom[36146] = 16'hffff;
  rom[36147] = 16'hffff;
  rom[36148] = 16'hffff;
  rom[36149] = 16'hffff;
  rom[36150] = 16'hffff;
  rom[36151] = 16'hffff;
  rom[36152] = 16'hffff;
  rom[36153] = 16'hffff;
  rom[36154] = 16'hffff;
  rom[36155] = 16'hffff;
  rom[36156] = 16'hffff;
  rom[36157] = 16'hffff;
  rom[36158] = 16'hffff;
  rom[36159] = 16'hffff;
  rom[36160] = 16'hffff;
  rom[36161] = 16'hffff;
  rom[36162] = 16'hffff;
  rom[36163] = 16'hffff;
  rom[36164] = 16'hffff;
  rom[36165] = 16'hffff;
  rom[36166] = 16'hffff;
  rom[36167] = 16'hffff;
  rom[36168] = 16'hffff;
  rom[36169] = 16'hffff;
  rom[36170] = 16'hffff;
  rom[36171] = 16'hffff;
  rom[36172] = 16'hffff;
  rom[36173] = 16'hffff;
  rom[36174] = 16'hffff;
  rom[36175] = 16'hffff;
  rom[36176] = 16'hffff;
  rom[36177] = 16'hffff;
  rom[36178] = 16'hffff;
  rom[36179] = 16'hffff;
  rom[36180] = 16'hffff;
  rom[36181] = 16'hffff;
  rom[36182] = 16'hffff;
  rom[36183] = 16'hffff;
  rom[36184] = 16'hffff;
  rom[36185] = 16'hffff;
  rom[36186] = 16'hffff;
  rom[36187] = 16'hffff;
  rom[36188] = 16'hffff;
  rom[36189] = 16'hffff;
  rom[36190] = 16'hffff;
  rom[36191] = 16'hffff;
  rom[36192] = 16'hffff;
  rom[36193] = 16'hffff;
  rom[36194] = 16'hffff;
  rom[36195] = 16'hffff;
  rom[36196] = 16'hffff;
  rom[36197] = 16'hffff;
  rom[36198] = 16'hffff;
  rom[36199] = 16'hffff;
  rom[36200] = 16'hffff;
  rom[36201] = 16'hffff;
  rom[36202] = 16'hffff;
  rom[36203] = 16'hffff;
  rom[36204] = 16'hffff;
  rom[36205] = 16'hffff;
  rom[36206] = 16'hffff;
  rom[36207] = 16'hffff;
  rom[36208] = 16'hffff;
  rom[36209] = 16'hffff;
  rom[36210] = 16'hffff;
  rom[36211] = 16'hffff;
  rom[36212] = 16'hffff;
  rom[36213] = 16'hffff;
  rom[36214] = 16'hffff;
  rom[36215] = 16'hffff;
  rom[36216] = 16'hffff;
  rom[36217] = 16'hffff;
  rom[36218] = 16'hffff;
  rom[36219] = 16'hffff;
  rom[36220] = 16'hffff;
  rom[36221] = 16'hffff;
  rom[36222] = 16'hffff;
  rom[36223] = 16'hffff;
  rom[36224] = 16'hffff;
  rom[36225] = 16'hffff;
  rom[36226] = 16'hffff;
  rom[36227] = 16'hffff;
  rom[36228] = 16'hffff;
  rom[36229] = 16'hffff;
  rom[36230] = 16'hffff;
  rom[36231] = 16'hffff;
  rom[36232] = 16'hffff;
  rom[36233] = 16'hffff;
  rom[36234] = 16'hffff;
  rom[36235] = 16'hffff;
  rom[36236] = 16'hffff;
  rom[36237] = 16'hffff;
  rom[36238] = 16'hffff;
  rom[36239] = 16'hffff;
  rom[36240] = 16'hffff;
  rom[36241] = 16'hffff;
  rom[36242] = 16'hffff;
  rom[36243] = 16'hffff;
  rom[36244] = 16'hffff;
  rom[36245] = 16'hffff;
  rom[36246] = 16'hffff;
  rom[36247] = 16'hffff;
  rom[36248] = 16'hffff;
  rom[36249] = 16'hffff;
  rom[36250] = 16'hffff;
  rom[36251] = 16'hffff;
  rom[36252] = 16'hffff;
  rom[36253] = 16'hffff;
  rom[36254] = 16'hffff;
  rom[36255] = 16'hffff;
  rom[36256] = 16'hffff;
  rom[36257] = 16'hffff;
  rom[36258] = 16'hffff;
  rom[36259] = 16'hffff;
  rom[36260] = 16'hffff;
  rom[36261] = 16'hffff;
  rom[36262] = 16'hffff;
  rom[36263] = 16'hffff;
  rom[36264] = 16'hffff;
  rom[36265] = 16'hffff;
  rom[36266] = 16'hffff;
  rom[36267] = 16'hffff;
  rom[36268] = 16'hffff;
  rom[36269] = 16'hffff;
  rom[36270] = 16'hffff;
  rom[36271] = 16'hffff;
  rom[36272] = 16'hffff;
  rom[36273] = 16'hffdf;
  rom[36274] = 16'hffde;
  rom[36275] = 16'h7387;
  rom[36276] = 16'hb548;
  rom[36277] = 16'hf74c;
  rom[36278] = 16'hff29;
  rom[36279] = 16'hf709;
  rom[36280] = 16'hff2a;
  rom[36281] = 16'hff28;
  rom[36282] = 16'hff49;
  rom[36283] = 16'hff29;
  rom[36284] = 16'hff29;
  rom[36285] = 16'hff28;
  rom[36286] = 16'hff28;
  rom[36287] = 16'hff28;
  rom[36288] = 16'hff29;
  rom[36289] = 16'hff29;
  rom[36290] = 16'hff29;
  rom[36291] = 16'hf728;
  rom[36292] = 16'hff2a;
  rom[36293] = 16'hff29;
  rom[36294] = 16'hff29;
  rom[36295] = 16'hff28;
  rom[36296] = 16'hff29;
  rom[36297] = 16'hff28;
  rom[36298] = 16'hff09;
  rom[36299] = 16'hff2d;
  rom[36300] = 16'h93a6;
  rom[36301] = 16'h7ac5;
  rom[36302] = 16'h9ba9;
  rom[36303] = 16'h8b68;
  rom[36304] = 16'h72c5;
  rom[36305] = 16'h6aa5;
  rom[36306] = 16'h8ba9;
  rom[36307] = 16'h8be9;
  rom[36308] = 16'h7b68;
  rom[36309] = 16'h8c6c;
  rom[36310] = 16'hdeb7;
  rom[36311] = 16'hffdc;
  rom[36312] = 16'hfffe;
  rom[36313] = 16'hffff;
  rom[36314] = 16'hffdf;
  rom[36315] = 16'hffbe;
  rom[36316] = 16'hffff;
  rom[36317] = 16'hffdf;
  rom[36318] = 16'hffff;
  rom[36319] = 16'hffff;
  rom[36320] = 16'hffff;
  rom[36321] = 16'hffff;
  rom[36322] = 16'hffff;
  rom[36323] = 16'hffff;
  rom[36324] = 16'hffff;
  rom[36325] = 16'hffff;
  rom[36326] = 16'hffff;
  rom[36327] = 16'hffff;
  rom[36328] = 16'hffff;
  rom[36329] = 16'hffff;
  rom[36330] = 16'hffff;
  rom[36331] = 16'hffff;
  rom[36332] = 16'hffff;
  rom[36333] = 16'hffff;
  rom[36334] = 16'hffff;
  rom[36335] = 16'hffff;
  rom[36336] = 16'hffff;
  rom[36337] = 16'hffff;
  rom[36338] = 16'hffff;
  rom[36339] = 16'hffff;
  rom[36340] = 16'hffff;
  rom[36341] = 16'hffff;
  rom[36342] = 16'hffff;
  rom[36343] = 16'hffff;
  rom[36344] = 16'hffff;
  rom[36345] = 16'hffff;
  rom[36346] = 16'hffff;
  rom[36347] = 16'hffff;
  rom[36348] = 16'hffff;
  rom[36349] = 16'hffff;
  rom[36350] = 16'hffff;
  rom[36351] = 16'hffff;
  rom[36352] = 16'hffff;
  rom[36353] = 16'hffff;
  rom[36354] = 16'hffff;
  rom[36355] = 16'hffff;
  rom[36356] = 16'hffff;
  rom[36357] = 16'hffff;
  rom[36358] = 16'hffff;
  rom[36359] = 16'hffff;
  rom[36360] = 16'hffff;
  rom[36361] = 16'hffff;
  rom[36362] = 16'hffff;
  rom[36363] = 16'hffff;
  rom[36364] = 16'hffff;
  rom[36365] = 16'hffff;
  rom[36366] = 16'hffff;
  rom[36367] = 16'hffff;
  rom[36368] = 16'hffff;
  rom[36369] = 16'hffff;
  rom[36370] = 16'hffff;
  rom[36371] = 16'hffff;
  rom[36372] = 16'hffff;
  rom[36373] = 16'hffff;
  rom[36374] = 16'hffff;
  rom[36375] = 16'hffff;
  rom[36376] = 16'hffff;
  rom[36377] = 16'hffff;
  rom[36378] = 16'hffff;
  rom[36379] = 16'hffff;
  rom[36380] = 16'hffff;
  rom[36381] = 16'hffff;
  rom[36382] = 16'hffff;
  rom[36383] = 16'hffff;
  rom[36384] = 16'hffff;
  rom[36385] = 16'hffff;
  rom[36386] = 16'hffff;
  rom[36387] = 16'hffff;
  rom[36388] = 16'hffff;
  rom[36389] = 16'hffff;
  rom[36390] = 16'hffff;
  rom[36391] = 16'hffff;
  rom[36392] = 16'hffff;
  rom[36393] = 16'hffff;
  rom[36394] = 16'hffff;
  rom[36395] = 16'hffff;
  rom[36396] = 16'hffff;
  rom[36397] = 16'hffff;
  rom[36398] = 16'hffff;
  rom[36399] = 16'hffff;
  rom[36400] = 16'hffff;
  rom[36401] = 16'hffff;
  rom[36402] = 16'hffff;
  rom[36403] = 16'hffff;
  rom[36404] = 16'hffff;
  rom[36405] = 16'hffff;
  rom[36406] = 16'hffff;
  rom[36407] = 16'hffff;
  rom[36408] = 16'hffff;
  rom[36409] = 16'hffff;
  rom[36410] = 16'hffff;
  rom[36411] = 16'hffff;
  rom[36412] = 16'hffff;
  rom[36413] = 16'hffff;
  rom[36414] = 16'hffff;
  rom[36415] = 16'hffff;
  rom[36416] = 16'hffff;
  rom[36417] = 16'hffff;
  rom[36418] = 16'hffff;
  rom[36419] = 16'hffff;
  rom[36420] = 16'hffff;
  rom[36421] = 16'hffff;
  rom[36422] = 16'hffff;
  rom[36423] = 16'hffff;
  rom[36424] = 16'hffff;
  rom[36425] = 16'hffff;
  rom[36426] = 16'hffff;
  rom[36427] = 16'hffff;
  rom[36428] = 16'hffff;
  rom[36429] = 16'hffff;
  rom[36430] = 16'hffff;
  rom[36431] = 16'hffff;
  rom[36432] = 16'hffff;
  rom[36433] = 16'hffff;
  rom[36434] = 16'hffff;
  rom[36435] = 16'hffff;
  rom[36436] = 16'hffff;
  rom[36437] = 16'hffff;
  rom[36438] = 16'hffff;
  rom[36439] = 16'hffff;
  rom[36440] = 16'hffff;
  rom[36441] = 16'hffff;
  rom[36442] = 16'hffff;
  rom[36443] = 16'hffff;
  rom[36444] = 16'hffff;
  rom[36445] = 16'hffff;
  rom[36446] = 16'hffff;
  rom[36447] = 16'hffff;
  rom[36448] = 16'hffff;
  rom[36449] = 16'hffff;
  rom[36450] = 16'hffff;
  rom[36451] = 16'hffff;
  rom[36452] = 16'hffff;
  rom[36453] = 16'hffff;
  rom[36454] = 16'hffff;
  rom[36455] = 16'hffff;
  rom[36456] = 16'hffff;
  rom[36457] = 16'hffff;
  rom[36458] = 16'hffff;
  rom[36459] = 16'hffff;
  rom[36460] = 16'hffff;
  rom[36461] = 16'hffff;
  rom[36462] = 16'hffff;
  rom[36463] = 16'hffff;
  rom[36464] = 16'hffff;
  rom[36465] = 16'hffff;
  rom[36466] = 16'hffff;
  rom[36467] = 16'hffff;
  rom[36468] = 16'hffff;
  rom[36469] = 16'hffff;
  rom[36470] = 16'hffff;
  rom[36471] = 16'hffff;
  rom[36472] = 16'hffff;
  rom[36473] = 16'hffdf;
  rom[36474] = 16'hffff;
  rom[36475] = 16'ha4ef;
  rom[36476] = 16'h7b84;
  rom[36477] = 16'heeec;
  rom[36478] = 16'hf72a;
  rom[36479] = 16'hff0a;
  rom[36480] = 16'hf709;
  rom[36481] = 16'hff28;
  rom[36482] = 16'hf708;
  rom[36483] = 16'hf709;
  rom[36484] = 16'hff09;
  rom[36485] = 16'hff29;
  rom[36486] = 16'hf708;
  rom[36487] = 16'hff28;
  rom[36488] = 16'hff08;
  rom[36489] = 16'hff29;
  rom[36490] = 16'hf708;
  rom[36491] = 16'hf749;
  rom[36492] = 16'hff09;
  rom[36493] = 16'hff29;
  rom[36494] = 16'hf708;
  rom[36495] = 16'hff28;
  rom[36496] = 16'hff08;
  rom[36497] = 16'hff29;
  rom[36498] = 16'hff29;
  rom[36499] = 16'hf70c;
  rom[36500] = 16'h9bc7;
  rom[36501] = 16'h8b6a;
  rom[36502] = 16'hde36;
  rom[36503] = 16'hf6f9;
  rom[36504] = 16'heed9;
  rom[36505] = 16'heefa;
  rom[36506] = 16'heef9;
  rom[36507] = 16'hef3a;
  rom[36508] = 16'hff9c;
  rom[36509] = 16'hfffe;
  rom[36510] = 16'hfffe;
  rom[36511] = 16'hffff;
  rom[36512] = 16'hffdf;
  rom[36513] = 16'hffff;
  rom[36514] = 16'hffff;
  rom[36515] = 16'hffff;
  rom[36516] = 16'hffff;
  rom[36517] = 16'hffff;
  rom[36518] = 16'hffff;
  rom[36519] = 16'hffff;
  rom[36520] = 16'hffff;
  rom[36521] = 16'hffff;
  rom[36522] = 16'hffff;
  rom[36523] = 16'hffff;
  rom[36524] = 16'hffff;
  rom[36525] = 16'hffff;
  rom[36526] = 16'hffff;
  rom[36527] = 16'hffff;
  rom[36528] = 16'hffff;
  rom[36529] = 16'hffff;
  rom[36530] = 16'hffff;
  rom[36531] = 16'hffff;
  rom[36532] = 16'hffff;
  rom[36533] = 16'hffff;
  rom[36534] = 16'hffff;
  rom[36535] = 16'hffff;
  rom[36536] = 16'hffff;
  rom[36537] = 16'hffff;
  rom[36538] = 16'hffff;
  rom[36539] = 16'hffff;
  rom[36540] = 16'hffff;
  rom[36541] = 16'hffff;
  rom[36542] = 16'hffff;
  rom[36543] = 16'hffff;
  rom[36544] = 16'hffff;
  rom[36545] = 16'hffff;
  rom[36546] = 16'hffff;
  rom[36547] = 16'hffff;
  rom[36548] = 16'hffff;
  rom[36549] = 16'hffff;
  rom[36550] = 16'hffff;
  rom[36551] = 16'hffff;
  rom[36552] = 16'hffff;
  rom[36553] = 16'hffff;
  rom[36554] = 16'hffff;
  rom[36555] = 16'hffff;
  rom[36556] = 16'hffff;
  rom[36557] = 16'hffff;
  rom[36558] = 16'hffff;
  rom[36559] = 16'hffff;
  rom[36560] = 16'hffff;
  rom[36561] = 16'hffff;
  rom[36562] = 16'hffff;
  rom[36563] = 16'hffff;
  rom[36564] = 16'hffff;
  rom[36565] = 16'hffff;
  rom[36566] = 16'hffff;
  rom[36567] = 16'hffff;
  rom[36568] = 16'hffff;
  rom[36569] = 16'hffff;
  rom[36570] = 16'hffff;
  rom[36571] = 16'hffff;
  rom[36572] = 16'hffff;
  rom[36573] = 16'hffff;
  rom[36574] = 16'hffff;
  rom[36575] = 16'hffff;
  rom[36576] = 16'hffff;
  rom[36577] = 16'hffff;
  rom[36578] = 16'hffff;
  rom[36579] = 16'hffff;
  rom[36580] = 16'hffff;
  rom[36581] = 16'hffff;
  rom[36582] = 16'hffff;
  rom[36583] = 16'hffff;
  rom[36584] = 16'hffff;
  rom[36585] = 16'hffff;
  rom[36586] = 16'hffff;
  rom[36587] = 16'hffff;
  rom[36588] = 16'hffff;
  rom[36589] = 16'hffff;
  rom[36590] = 16'hffff;
  rom[36591] = 16'hffff;
  rom[36592] = 16'hffff;
  rom[36593] = 16'hffff;
  rom[36594] = 16'hffff;
  rom[36595] = 16'hffff;
  rom[36596] = 16'hffff;
  rom[36597] = 16'hffff;
  rom[36598] = 16'hffff;
  rom[36599] = 16'hffff;
  rom[36600] = 16'hffff;
  rom[36601] = 16'hffff;
  rom[36602] = 16'hffff;
  rom[36603] = 16'hffff;
  rom[36604] = 16'hffff;
  rom[36605] = 16'hffff;
  rom[36606] = 16'hffff;
  rom[36607] = 16'hffff;
  rom[36608] = 16'hffff;
  rom[36609] = 16'hffff;
  rom[36610] = 16'hffff;
  rom[36611] = 16'hffff;
  rom[36612] = 16'hffff;
  rom[36613] = 16'hffff;
  rom[36614] = 16'hffff;
  rom[36615] = 16'hffff;
  rom[36616] = 16'hffff;
  rom[36617] = 16'hffff;
  rom[36618] = 16'hffff;
  rom[36619] = 16'hffff;
  rom[36620] = 16'hffff;
  rom[36621] = 16'hffff;
  rom[36622] = 16'hffff;
  rom[36623] = 16'hffff;
  rom[36624] = 16'hffff;
  rom[36625] = 16'hffff;
  rom[36626] = 16'hffff;
  rom[36627] = 16'hffff;
  rom[36628] = 16'hffff;
  rom[36629] = 16'hffff;
  rom[36630] = 16'hffff;
  rom[36631] = 16'hffff;
  rom[36632] = 16'hffff;
  rom[36633] = 16'hffff;
  rom[36634] = 16'hffff;
  rom[36635] = 16'hffff;
  rom[36636] = 16'hffff;
  rom[36637] = 16'hffff;
  rom[36638] = 16'hffff;
  rom[36639] = 16'hffff;
  rom[36640] = 16'hffff;
  rom[36641] = 16'hffff;
  rom[36642] = 16'hffff;
  rom[36643] = 16'hffff;
  rom[36644] = 16'hffff;
  rom[36645] = 16'hffff;
  rom[36646] = 16'hffff;
  rom[36647] = 16'hffff;
  rom[36648] = 16'hffff;
  rom[36649] = 16'hffff;
  rom[36650] = 16'hffff;
  rom[36651] = 16'hffff;
  rom[36652] = 16'hffff;
  rom[36653] = 16'hffff;
  rom[36654] = 16'hffff;
  rom[36655] = 16'hffff;
  rom[36656] = 16'hffff;
  rom[36657] = 16'hffff;
  rom[36658] = 16'hffff;
  rom[36659] = 16'hffff;
  rom[36660] = 16'hffff;
  rom[36661] = 16'hffff;
  rom[36662] = 16'hffff;
  rom[36663] = 16'hffff;
  rom[36664] = 16'hffff;
  rom[36665] = 16'hffff;
  rom[36666] = 16'hffff;
  rom[36667] = 16'hffff;
  rom[36668] = 16'hffff;
  rom[36669] = 16'hffff;
  rom[36670] = 16'hffff;
  rom[36671] = 16'hffff;
  rom[36672] = 16'hffff;
  rom[36673] = 16'hffff;
  rom[36674] = 16'hffdf;
  rom[36675] = 16'hbdd5;
  rom[36676] = 16'h5a61;
  rom[36677] = 16'he68d;
  rom[36678] = 16'hff2b;
  rom[36679] = 16'hff0a;
  rom[36680] = 16'hff0a;
  rom[36681] = 16'hff28;
  rom[36682] = 16'hff49;
  rom[36683] = 16'hf709;
  rom[36684] = 16'hff2a;
  rom[36685] = 16'hff29;
  rom[36686] = 16'hff29;
  rom[36687] = 16'hff28;
  rom[36688] = 16'hff29;
  rom[36689] = 16'hff29;
  rom[36690] = 16'hff29;
  rom[36691] = 16'hff28;
  rom[36692] = 16'hff2a;
  rom[36693] = 16'hff29;
  rom[36694] = 16'hff29;
  rom[36695] = 16'hff28;
  rom[36696] = 16'hff29;
  rom[36697] = 16'hf708;
  rom[36698] = 16'hff2a;
  rom[36699] = 16'hf70c;
  rom[36700] = 16'h8ba8;
  rom[36701] = 16'h9c2d;
  rom[36702] = 16'hffde;
  rom[36703] = 16'hfffe;
  rom[36704] = 16'hffff;
  rom[36705] = 16'hffff;
  rom[36706] = 16'hffff;
  rom[36707] = 16'hffff;
  rom[36708] = 16'hffff;
  rom[36709] = 16'hffff;
  rom[36710] = 16'hffff;
  rom[36711] = 16'hffff;
  rom[36712] = 16'hffff;
  rom[36713] = 16'hffff;
  rom[36714] = 16'hffff;
  rom[36715] = 16'hffff;
  rom[36716] = 16'hffff;
  rom[36717] = 16'hffff;
  rom[36718] = 16'hffff;
  rom[36719] = 16'hffff;
  rom[36720] = 16'hffff;
  rom[36721] = 16'hffff;
  rom[36722] = 16'hffff;
  rom[36723] = 16'hffff;
  rom[36724] = 16'hffff;
  rom[36725] = 16'hffff;
  rom[36726] = 16'hffff;
  rom[36727] = 16'hffff;
  rom[36728] = 16'hffff;
  rom[36729] = 16'hffff;
  rom[36730] = 16'hffff;
  rom[36731] = 16'hffff;
  rom[36732] = 16'hffff;
  rom[36733] = 16'hffff;
  rom[36734] = 16'hffff;
  rom[36735] = 16'hffff;
  rom[36736] = 16'hffff;
  rom[36737] = 16'hffff;
  rom[36738] = 16'hffff;
  rom[36739] = 16'hffff;
  rom[36740] = 16'hffff;
  rom[36741] = 16'hffff;
  rom[36742] = 16'hffff;
  rom[36743] = 16'hffff;
  rom[36744] = 16'hffff;
  rom[36745] = 16'hffff;
  rom[36746] = 16'hffff;
  rom[36747] = 16'hffff;
  rom[36748] = 16'hffff;
  rom[36749] = 16'hffff;
  rom[36750] = 16'hffff;
  rom[36751] = 16'hffff;
  rom[36752] = 16'hffff;
  rom[36753] = 16'hffff;
  rom[36754] = 16'hffff;
  rom[36755] = 16'hffff;
  rom[36756] = 16'hffff;
  rom[36757] = 16'hffff;
  rom[36758] = 16'hffff;
  rom[36759] = 16'hffff;
  rom[36760] = 16'hffff;
  rom[36761] = 16'hffff;
  rom[36762] = 16'hffff;
  rom[36763] = 16'hffff;
  rom[36764] = 16'hffff;
  rom[36765] = 16'hffff;
  rom[36766] = 16'hffff;
  rom[36767] = 16'hffff;
  rom[36768] = 16'hffff;
  rom[36769] = 16'hffff;
  rom[36770] = 16'hffff;
  rom[36771] = 16'hffff;
  rom[36772] = 16'hffff;
  rom[36773] = 16'hffff;
  rom[36774] = 16'hffff;
  rom[36775] = 16'hffff;
  rom[36776] = 16'hffff;
  rom[36777] = 16'hffff;
  rom[36778] = 16'hffff;
  rom[36779] = 16'hffff;
  rom[36780] = 16'hffff;
  rom[36781] = 16'hffff;
  rom[36782] = 16'hffff;
  rom[36783] = 16'hffff;
  rom[36784] = 16'hffff;
  rom[36785] = 16'hffff;
  rom[36786] = 16'hffff;
  rom[36787] = 16'hffff;
  rom[36788] = 16'hffff;
  rom[36789] = 16'hffff;
  rom[36790] = 16'hffff;
  rom[36791] = 16'hffff;
  rom[36792] = 16'hffff;
  rom[36793] = 16'hffff;
  rom[36794] = 16'hffff;
  rom[36795] = 16'hffff;
  rom[36796] = 16'hffff;
  rom[36797] = 16'hffff;
  rom[36798] = 16'hffff;
  rom[36799] = 16'hffff;
  rom[36800] = 16'hffff;
  rom[36801] = 16'hffff;
  rom[36802] = 16'hffff;
  rom[36803] = 16'hffff;
  rom[36804] = 16'hffff;
  rom[36805] = 16'hffff;
  rom[36806] = 16'hffff;
  rom[36807] = 16'hffff;
  rom[36808] = 16'hffff;
  rom[36809] = 16'hffff;
  rom[36810] = 16'hffff;
  rom[36811] = 16'hffff;
  rom[36812] = 16'hffff;
  rom[36813] = 16'hffff;
  rom[36814] = 16'hffff;
  rom[36815] = 16'hffff;
  rom[36816] = 16'hffff;
  rom[36817] = 16'hffff;
  rom[36818] = 16'hffff;
  rom[36819] = 16'hffff;
  rom[36820] = 16'hffff;
  rom[36821] = 16'hffff;
  rom[36822] = 16'hffff;
  rom[36823] = 16'hffff;
  rom[36824] = 16'hffff;
  rom[36825] = 16'hffff;
  rom[36826] = 16'hffff;
  rom[36827] = 16'hffff;
  rom[36828] = 16'hffff;
  rom[36829] = 16'hffff;
  rom[36830] = 16'hffff;
  rom[36831] = 16'hffff;
  rom[36832] = 16'hffff;
  rom[36833] = 16'hffff;
  rom[36834] = 16'hffff;
  rom[36835] = 16'hffff;
  rom[36836] = 16'hffff;
  rom[36837] = 16'hffff;
  rom[36838] = 16'hffff;
  rom[36839] = 16'hffff;
  rom[36840] = 16'hffff;
  rom[36841] = 16'hffff;
  rom[36842] = 16'hffff;
  rom[36843] = 16'hffff;
  rom[36844] = 16'hffff;
  rom[36845] = 16'hffff;
  rom[36846] = 16'hffff;
  rom[36847] = 16'hffff;
  rom[36848] = 16'hffff;
  rom[36849] = 16'hffff;
  rom[36850] = 16'hffff;
  rom[36851] = 16'hffff;
  rom[36852] = 16'hffff;
  rom[36853] = 16'hffff;
  rom[36854] = 16'hffff;
  rom[36855] = 16'hffff;
  rom[36856] = 16'hffff;
  rom[36857] = 16'hffff;
  rom[36858] = 16'hffff;
  rom[36859] = 16'hffff;
  rom[36860] = 16'hffff;
  rom[36861] = 16'hffff;
  rom[36862] = 16'hffff;
  rom[36863] = 16'hffff;
  rom[36864] = 16'hffff;
  rom[36865] = 16'hffff;
  rom[36866] = 16'hffff;
  rom[36867] = 16'hffff;
  rom[36868] = 16'hffff;
  rom[36869] = 16'hffff;
  rom[36870] = 16'hffff;
  rom[36871] = 16'hffff;
  rom[36872] = 16'hfffe;
  rom[36873] = 16'hffff;
  rom[36874] = 16'hffff;
  rom[36875] = 16'he6db;
  rom[36876] = 16'h49e2;
  rom[36877] = 16'hbd8a;
  rom[36878] = 16'hf72c;
  rom[36879] = 16'hff0a;
  rom[36880] = 16'hff09;
  rom[36881] = 16'hff08;
  rom[36882] = 16'hff28;
  rom[36883] = 16'hff29;
  rom[36884] = 16'hf709;
  rom[36885] = 16'hff29;
  rom[36886] = 16'hff08;
  rom[36887] = 16'hff28;
  rom[36888] = 16'hf708;
  rom[36889] = 16'hff29;
  rom[36890] = 16'hff08;
  rom[36891] = 16'hff29;
  rom[36892] = 16'hf709;
  rom[36893] = 16'hff29;
  rom[36894] = 16'hff08;
  rom[36895] = 16'hff28;
  rom[36896] = 16'hff08;
  rom[36897] = 16'hff28;
  rom[36898] = 16'hff4a;
  rom[36899] = 16'hf70c;
  rom[36900] = 16'h7b65;
  rom[36901] = 16'h944e;
  rom[36902] = 16'hffbd;
  rom[36903] = 16'hffff;
  rom[36904] = 16'hffff;
  rom[36905] = 16'hffff;
  rom[36906] = 16'hffff;
  rom[36907] = 16'hffff;
  rom[36908] = 16'hffff;
  rom[36909] = 16'hffff;
  rom[36910] = 16'hffff;
  rom[36911] = 16'hffff;
  rom[36912] = 16'hffff;
  rom[36913] = 16'hffff;
  rom[36914] = 16'hffff;
  rom[36915] = 16'hffff;
  rom[36916] = 16'hffff;
  rom[36917] = 16'hffff;
  rom[36918] = 16'hffff;
  rom[36919] = 16'hffff;
  rom[36920] = 16'hffff;
  rom[36921] = 16'hffff;
  rom[36922] = 16'hffff;
  rom[36923] = 16'hffff;
  rom[36924] = 16'hffff;
  rom[36925] = 16'hffff;
  rom[36926] = 16'hffff;
  rom[36927] = 16'hffff;
  rom[36928] = 16'hffff;
  rom[36929] = 16'hffff;
  rom[36930] = 16'hffff;
  rom[36931] = 16'hffff;
  rom[36932] = 16'hffff;
  rom[36933] = 16'hffff;
  rom[36934] = 16'hffff;
  rom[36935] = 16'hffff;
  rom[36936] = 16'hffff;
  rom[36937] = 16'hffff;
  rom[36938] = 16'hffff;
  rom[36939] = 16'hffff;
  rom[36940] = 16'hffff;
  rom[36941] = 16'hffff;
  rom[36942] = 16'hffff;
  rom[36943] = 16'hffff;
  rom[36944] = 16'hffff;
  rom[36945] = 16'hffff;
  rom[36946] = 16'hffff;
  rom[36947] = 16'hffff;
  rom[36948] = 16'hffff;
  rom[36949] = 16'hffff;
  rom[36950] = 16'hffff;
  rom[36951] = 16'hffff;
  rom[36952] = 16'hffff;
  rom[36953] = 16'hffff;
  rom[36954] = 16'hffff;
  rom[36955] = 16'hffff;
  rom[36956] = 16'hffff;
  rom[36957] = 16'hffff;
  rom[36958] = 16'hffff;
  rom[36959] = 16'hffff;
  rom[36960] = 16'hffff;
  rom[36961] = 16'hffff;
  rom[36962] = 16'hffff;
  rom[36963] = 16'hffff;
  rom[36964] = 16'hffff;
  rom[36965] = 16'hffff;
  rom[36966] = 16'hffff;
  rom[36967] = 16'hffff;
  rom[36968] = 16'hffff;
  rom[36969] = 16'hffff;
  rom[36970] = 16'hffff;
  rom[36971] = 16'hffff;
  rom[36972] = 16'hffff;
  rom[36973] = 16'hffff;
  rom[36974] = 16'hffff;
  rom[36975] = 16'hffff;
  rom[36976] = 16'hffff;
  rom[36977] = 16'hffff;
  rom[36978] = 16'hffff;
  rom[36979] = 16'hffff;
  rom[36980] = 16'hffff;
  rom[36981] = 16'hffff;
  rom[36982] = 16'hffff;
  rom[36983] = 16'hffff;
  rom[36984] = 16'hffff;
  rom[36985] = 16'hffff;
  rom[36986] = 16'hffff;
  rom[36987] = 16'hffff;
  rom[36988] = 16'hffff;
  rom[36989] = 16'hffff;
  rom[36990] = 16'hffff;
  rom[36991] = 16'hffff;
  rom[36992] = 16'hffff;
  rom[36993] = 16'hffff;
  rom[36994] = 16'hffff;
  rom[36995] = 16'hffff;
  rom[36996] = 16'hffff;
  rom[36997] = 16'hffff;
  rom[36998] = 16'hffff;
  rom[36999] = 16'hffff;
  rom[37000] = 16'hffff;
  rom[37001] = 16'hffff;
  rom[37002] = 16'hffff;
  rom[37003] = 16'hffff;
  rom[37004] = 16'hffff;
  rom[37005] = 16'hffff;
  rom[37006] = 16'hffff;
  rom[37007] = 16'hffff;
  rom[37008] = 16'hffff;
  rom[37009] = 16'hffff;
  rom[37010] = 16'hffff;
  rom[37011] = 16'hffff;
  rom[37012] = 16'hffff;
  rom[37013] = 16'hffff;
  rom[37014] = 16'hffff;
  rom[37015] = 16'hffff;
  rom[37016] = 16'hffff;
  rom[37017] = 16'hffff;
  rom[37018] = 16'hffff;
  rom[37019] = 16'hffff;
  rom[37020] = 16'hffff;
  rom[37021] = 16'hffff;
  rom[37022] = 16'hffff;
  rom[37023] = 16'hffff;
  rom[37024] = 16'hffff;
  rom[37025] = 16'hffff;
  rom[37026] = 16'hffff;
  rom[37027] = 16'hffff;
  rom[37028] = 16'hffff;
  rom[37029] = 16'hffff;
  rom[37030] = 16'hffff;
  rom[37031] = 16'hffff;
  rom[37032] = 16'hffff;
  rom[37033] = 16'hffff;
  rom[37034] = 16'hffff;
  rom[37035] = 16'hffff;
  rom[37036] = 16'hffff;
  rom[37037] = 16'hffff;
  rom[37038] = 16'hffff;
  rom[37039] = 16'hffff;
  rom[37040] = 16'hffff;
  rom[37041] = 16'hffff;
  rom[37042] = 16'hffff;
  rom[37043] = 16'hffff;
  rom[37044] = 16'hffff;
  rom[37045] = 16'hffff;
  rom[37046] = 16'hffff;
  rom[37047] = 16'hffff;
  rom[37048] = 16'hffff;
  rom[37049] = 16'hffff;
  rom[37050] = 16'hffff;
  rom[37051] = 16'hffff;
  rom[37052] = 16'hffff;
  rom[37053] = 16'hffff;
  rom[37054] = 16'hffff;
  rom[37055] = 16'hffff;
  rom[37056] = 16'hffff;
  rom[37057] = 16'hffff;
  rom[37058] = 16'hffff;
  rom[37059] = 16'hffff;
  rom[37060] = 16'hffff;
  rom[37061] = 16'hffff;
  rom[37062] = 16'hffff;
  rom[37063] = 16'hffff;
  rom[37064] = 16'hffff;
  rom[37065] = 16'hffff;
  rom[37066] = 16'hffff;
  rom[37067] = 16'hffff;
  rom[37068] = 16'hffff;
  rom[37069] = 16'hffff;
  rom[37070] = 16'hffff;
  rom[37071] = 16'hffff;
  rom[37072] = 16'hffff;
  rom[37073] = 16'hffff;
  rom[37074] = 16'hffff;
  rom[37075] = 16'hffdf;
  rom[37076] = 16'h7348;
  rom[37077] = 16'h83e5;
  rom[37078] = 16'hff4d;
  rom[37079] = 16'hf6c9;
  rom[37080] = 16'hff2a;
  rom[37081] = 16'hff08;
  rom[37082] = 16'hff29;
  rom[37083] = 16'hff29;
  rom[37084] = 16'hff2a;
  rom[37085] = 16'hff29;
  rom[37086] = 16'hff29;
  rom[37087] = 16'hff28;
  rom[37088] = 16'hff49;
  rom[37089] = 16'hff28;
  rom[37090] = 16'hff29;
  rom[37091] = 16'hff28;
  rom[37092] = 16'hff2a;
  rom[37093] = 16'hff29;
  rom[37094] = 16'hff29;
  rom[37095] = 16'hff28;
  rom[37096] = 16'hff29;
  rom[37097] = 16'hff09;
  rom[37098] = 16'hff4a;
  rom[37099] = 16'hef0d;
  rom[37100] = 16'h7b45;
  rom[37101] = 16'ha4d0;
  rom[37102] = 16'hfffe;
  rom[37103] = 16'hffff;
  rom[37104] = 16'hffff;
  rom[37105] = 16'hffff;
  rom[37106] = 16'hffff;
  rom[37107] = 16'hffff;
  rom[37108] = 16'hffff;
  rom[37109] = 16'hffff;
  rom[37110] = 16'hffff;
  rom[37111] = 16'hffff;
  rom[37112] = 16'hffff;
  rom[37113] = 16'hffff;
  rom[37114] = 16'hffff;
  rom[37115] = 16'hffff;
  rom[37116] = 16'hffff;
  rom[37117] = 16'hffff;
  rom[37118] = 16'hffff;
  rom[37119] = 16'hffff;
  rom[37120] = 16'hffff;
  rom[37121] = 16'hffff;
  rom[37122] = 16'hffff;
  rom[37123] = 16'hffff;
  rom[37124] = 16'hffff;
  rom[37125] = 16'hffff;
  rom[37126] = 16'hffff;
  rom[37127] = 16'hffff;
  rom[37128] = 16'hffff;
  rom[37129] = 16'hffff;
  rom[37130] = 16'hffff;
  rom[37131] = 16'hffff;
  rom[37132] = 16'hffff;
  rom[37133] = 16'hffff;
  rom[37134] = 16'hffff;
  rom[37135] = 16'hffff;
  rom[37136] = 16'hffff;
  rom[37137] = 16'hffff;
  rom[37138] = 16'hffff;
  rom[37139] = 16'hffff;
  rom[37140] = 16'hffff;
  rom[37141] = 16'hffff;
  rom[37142] = 16'hffff;
  rom[37143] = 16'hffff;
  rom[37144] = 16'hffff;
  rom[37145] = 16'hffff;
  rom[37146] = 16'hffff;
  rom[37147] = 16'hffff;
  rom[37148] = 16'hffff;
  rom[37149] = 16'hffff;
  rom[37150] = 16'hffff;
  rom[37151] = 16'hffff;
  rom[37152] = 16'hffff;
  rom[37153] = 16'hffff;
  rom[37154] = 16'hffff;
  rom[37155] = 16'hffff;
  rom[37156] = 16'hffff;
  rom[37157] = 16'hffff;
  rom[37158] = 16'hffff;
  rom[37159] = 16'hffff;
  rom[37160] = 16'hffff;
  rom[37161] = 16'hffff;
  rom[37162] = 16'hffff;
  rom[37163] = 16'hffff;
  rom[37164] = 16'hffff;
  rom[37165] = 16'hffff;
  rom[37166] = 16'hffff;
  rom[37167] = 16'hffff;
  rom[37168] = 16'hffff;
  rom[37169] = 16'hffff;
  rom[37170] = 16'hffff;
  rom[37171] = 16'hffff;
  rom[37172] = 16'hffff;
  rom[37173] = 16'hffff;
  rom[37174] = 16'hffff;
  rom[37175] = 16'hffff;
  rom[37176] = 16'hffff;
  rom[37177] = 16'hffff;
  rom[37178] = 16'hffff;
  rom[37179] = 16'hffff;
  rom[37180] = 16'hffff;
  rom[37181] = 16'hffff;
  rom[37182] = 16'hffff;
  rom[37183] = 16'hffff;
  rom[37184] = 16'hffff;
  rom[37185] = 16'hffff;
  rom[37186] = 16'hffff;
  rom[37187] = 16'hffff;
  rom[37188] = 16'hffff;
  rom[37189] = 16'hffff;
  rom[37190] = 16'hffff;
  rom[37191] = 16'hffff;
  rom[37192] = 16'hffff;
  rom[37193] = 16'hffff;
  rom[37194] = 16'hffff;
  rom[37195] = 16'hffff;
  rom[37196] = 16'hffff;
  rom[37197] = 16'hffff;
  rom[37198] = 16'hffff;
  rom[37199] = 16'hffff;
  rom[37200] = 16'hffff;
  rom[37201] = 16'hffff;
  rom[37202] = 16'hffff;
  rom[37203] = 16'hffff;
  rom[37204] = 16'hffff;
  rom[37205] = 16'hffff;
  rom[37206] = 16'hffff;
  rom[37207] = 16'hffff;
  rom[37208] = 16'hffff;
  rom[37209] = 16'hffff;
  rom[37210] = 16'hffff;
  rom[37211] = 16'hffff;
  rom[37212] = 16'hffff;
  rom[37213] = 16'hffff;
  rom[37214] = 16'hffff;
  rom[37215] = 16'hffff;
  rom[37216] = 16'hffff;
  rom[37217] = 16'hffff;
  rom[37218] = 16'hffff;
  rom[37219] = 16'hffff;
  rom[37220] = 16'hffff;
  rom[37221] = 16'hffff;
  rom[37222] = 16'hffff;
  rom[37223] = 16'hffff;
  rom[37224] = 16'hffff;
  rom[37225] = 16'hffff;
  rom[37226] = 16'hffff;
  rom[37227] = 16'hffff;
  rom[37228] = 16'hffff;
  rom[37229] = 16'hffff;
  rom[37230] = 16'hffff;
  rom[37231] = 16'hffff;
  rom[37232] = 16'hffff;
  rom[37233] = 16'hffff;
  rom[37234] = 16'hffff;
  rom[37235] = 16'hffff;
  rom[37236] = 16'hffff;
  rom[37237] = 16'hffff;
  rom[37238] = 16'hffff;
  rom[37239] = 16'hffff;
  rom[37240] = 16'hffff;
  rom[37241] = 16'hffff;
  rom[37242] = 16'hffff;
  rom[37243] = 16'hffff;
  rom[37244] = 16'hffff;
  rom[37245] = 16'hffff;
  rom[37246] = 16'hffff;
  rom[37247] = 16'hffff;
  rom[37248] = 16'hffff;
  rom[37249] = 16'hffff;
  rom[37250] = 16'hffff;
  rom[37251] = 16'hffff;
  rom[37252] = 16'hffff;
  rom[37253] = 16'hffff;
  rom[37254] = 16'hffff;
  rom[37255] = 16'hffff;
  rom[37256] = 16'hffff;
  rom[37257] = 16'hffff;
  rom[37258] = 16'hffff;
  rom[37259] = 16'hffff;
  rom[37260] = 16'hffff;
  rom[37261] = 16'hffff;
  rom[37262] = 16'hffff;
  rom[37263] = 16'hffff;
  rom[37264] = 16'hffff;
  rom[37265] = 16'hffff;
  rom[37266] = 16'hffff;
  rom[37267] = 16'hffff;
  rom[37268] = 16'hffff;
  rom[37269] = 16'hffff;
  rom[37270] = 16'hffff;
  rom[37271] = 16'hffff;
  rom[37272] = 16'hffff;
  rom[37273] = 16'hffff;
  rom[37274] = 16'hffdf;
  rom[37275] = 16'hffdf;
  rom[37276] = 16'hb551;
  rom[37277] = 16'h62e3;
  rom[37278] = 16'he6cc;
  rom[37279] = 16'hf70a;
  rom[37280] = 16'hf709;
  rom[37281] = 16'hff49;
  rom[37282] = 16'hf728;
  rom[37283] = 16'hff29;
  rom[37284] = 16'hf708;
  rom[37285] = 16'hff29;
  rom[37286] = 16'hf708;
  rom[37287] = 16'hff28;
  rom[37288] = 16'hff28;
  rom[37289] = 16'hff28;
  rom[37290] = 16'hf708;
  rom[37291] = 16'hff29;
  rom[37292] = 16'hff09;
  rom[37293] = 16'hf729;
  rom[37294] = 16'hf708;
  rom[37295] = 16'hff28;
  rom[37296] = 16'hff09;
  rom[37297] = 16'hff29;
  rom[37298] = 16'hf709;
  rom[37299] = 16'hf74d;
  rom[37300] = 16'h6b05;
  rom[37301] = 16'hb532;
  rom[37302] = 16'hfffe;
  rom[37303] = 16'hffff;
  rom[37304] = 16'hffff;
  rom[37305] = 16'hffff;
  rom[37306] = 16'hffff;
  rom[37307] = 16'hffff;
  rom[37308] = 16'hffff;
  rom[37309] = 16'hffff;
  rom[37310] = 16'hffff;
  rom[37311] = 16'hffff;
  rom[37312] = 16'hffff;
  rom[37313] = 16'hffff;
  rom[37314] = 16'hffff;
  rom[37315] = 16'hffff;
  rom[37316] = 16'hffff;
  rom[37317] = 16'hffff;
  rom[37318] = 16'hffff;
  rom[37319] = 16'hffff;
  rom[37320] = 16'hffff;
  rom[37321] = 16'hffff;
  rom[37322] = 16'hffff;
  rom[37323] = 16'hffff;
  rom[37324] = 16'hffff;
  rom[37325] = 16'hffff;
  rom[37326] = 16'hffff;
  rom[37327] = 16'hffff;
  rom[37328] = 16'hffff;
  rom[37329] = 16'hffff;
  rom[37330] = 16'hffff;
  rom[37331] = 16'hffff;
  rom[37332] = 16'hffff;
  rom[37333] = 16'hffff;
  rom[37334] = 16'hffff;
  rom[37335] = 16'hffff;
  rom[37336] = 16'hffff;
  rom[37337] = 16'hffff;
  rom[37338] = 16'hffff;
  rom[37339] = 16'hffff;
  rom[37340] = 16'hffff;
  rom[37341] = 16'hffff;
  rom[37342] = 16'hffff;
  rom[37343] = 16'hffff;
  rom[37344] = 16'hffff;
  rom[37345] = 16'hffff;
  rom[37346] = 16'hffff;
  rom[37347] = 16'hffff;
  rom[37348] = 16'hffff;
  rom[37349] = 16'hffff;
  rom[37350] = 16'hffff;
  rom[37351] = 16'hffff;
  rom[37352] = 16'hffff;
  rom[37353] = 16'hffff;
  rom[37354] = 16'hffff;
  rom[37355] = 16'hffff;
  rom[37356] = 16'hffff;
  rom[37357] = 16'hffff;
  rom[37358] = 16'hffff;
  rom[37359] = 16'hffff;
  rom[37360] = 16'hffff;
  rom[37361] = 16'hffff;
  rom[37362] = 16'hffff;
  rom[37363] = 16'hffff;
  rom[37364] = 16'hffff;
  rom[37365] = 16'hffff;
  rom[37366] = 16'hffff;
  rom[37367] = 16'hffff;
  rom[37368] = 16'hffff;
  rom[37369] = 16'hffff;
  rom[37370] = 16'hffff;
  rom[37371] = 16'hffff;
  rom[37372] = 16'hffff;
  rom[37373] = 16'hffff;
  rom[37374] = 16'hffff;
  rom[37375] = 16'hffff;
  rom[37376] = 16'hffff;
  rom[37377] = 16'hffff;
  rom[37378] = 16'hffff;
  rom[37379] = 16'hffff;
  rom[37380] = 16'hffff;
  rom[37381] = 16'hffff;
  rom[37382] = 16'hffff;
  rom[37383] = 16'hffff;
  rom[37384] = 16'hffff;
  rom[37385] = 16'hffff;
  rom[37386] = 16'hffff;
  rom[37387] = 16'hffff;
  rom[37388] = 16'hffff;
  rom[37389] = 16'hffff;
  rom[37390] = 16'hffff;
  rom[37391] = 16'hffff;
  rom[37392] = 16'hffff;
  rom[37393] = 16'hffff;
  rom[37394] = 16'hffff;
  rom[37395] = 16'hffff;
  rom[37396] = 16'hffff;
  rom[37397] = 16'hffff;
  rom[37398] = 16'hffff;
  rom[37399] = 16'hffff;
  rom[37400] = 16'hffff;
  rom[37401] = 16'hffff;
  rom[37402] = 16'hffff;
  rom[37403] = 16'hffff;
  rom[37404] = 16'hffff;
  rom[37405] = 16'hffff;
  rom[37406] = 16'hffff;
  rom[37407] = 16'hffff;
  rom[37408] = 16'hffff;
  rom[37409] = 16'hffff;
  rom[37410] = 16'hffff;
  rom[37411] = 16'hffff;
  rom[37412] = 16'hffff;
  rom[37413] = 16'hffff;
  rom[37414] = 16'hffff;
  rom[37415] = 16'hffff;
  rom[37416] = 16'hffff;
  rom[37417] = 16'hffff;
  rom[37418] = 16'hffff;
  rom[37419] = 16'hffff;
  rom[37420] = 16'hffff;
  rom[37421] = 16'hffff;
  rom[37422] = 16'hffff;
  rom[37423] = 16'hffff;
  rom[37424] = 16'hffff;
  rom[37425] = 16'hffff;
  rom[37426] = 16'hffff;
  rom[37427] = 16'hffff;
  rom[37428] = 16'hffff;
  rom[37429] = 16'hffff;
  rom[37430] = 16'hffff;
  rom[37431] = 16'hffff;
  rom[37432] = 16'hffff;
  rom[37433] = 16'hffff;
  rom[37434] = 16'hffff;
  rom[37435] = 16'hffff;
  rom[37436] = 16'hffff;
  rom[37437] = 16'hffff;
  rom[37438] = 16'hffff;
  rom[37439] = 16'hffff;
  rom[37440] = 16'hffff;
  rom[37441] = 16'hffff;
  rom[37442] = 16'hffff;
  rom[37443] = 16'hffff;
  rom[37444] = 16'hffff;
  rom[37445] = 16'hffff;
  rom[37446] = 16'hffff;
  rom[37447] = 16'hffff;
  rom[37448] = 16'hffff;
  rom[37449] = 16'hffff;
  rom[37450] = 16'hffff;
  rom[37451] = 16'hffff;
  rom[37452] = 16'hffff;
  rom[37453] = 16'hffff;
  rom[37454] = 16'hffff;
  rom[37455] = 16'hffff;
  rom[37456] = 16'hffff;
  rom[37457] = 16'hffff;
  rom[37458] = 16'hffff;
  rom[37459] = 16'hffff;
  rom[37460] = 16'hffff;
  rom[37461] = 16'hffff;
  rom[37462] = 16'hffff;
  rom[37463] = 16'hffff;
  rom[37464] = 16'hffff;
  rom[37465] = 16'hffff;
  rom[37466] = 16'hffff;
  rom[37467] = 16'hffff;
  rom[37468] = 16'hffff;
  rom[37469] = 16'hffff;
  rom[37470] = 16'hffff;
  rom[37471] = 16'hffff;
  rom[37472] = 16'hffff;
  rom[37473] = 16'hffff;
  rom[37474] = 16'hffff;
  rom[37475] = 16'hffdf;
  rom[37476] = 16'hff9c;
  rom[37477] = 16'h5a82;
  rom[37478] = 16'hd62b;
  rom[37479] = 16'hf72c;
  rom[37480] = 16'hff2a;
  rom[37481] = 16'hff49;
  rom[37482] = 16'hff28;
  rom[37483] = 16'hf708;
  rom[37484] = 16'hff4a;
  rom[37485] = 16'hff29;
  rom[37486] = 16'hff29;
  rom[37487] = 16'hff28;
  rom[37488] = 16'hff49;
  rom[37489] = 16'hff28;
  rom[37490] = 16'hff29;
  rom[37491] = 16'hff28;
  rom[37492] = 16'hff2a;
  rom[37493] = 16'hf729;
  rom[37494] = 16'hff29;
  rom[37495] = 16'hff28;
  rom[37496] = 16'hff2a;
  rom[37497] = 16'hff29;
  rom[37498] = 16'hf709;
  rom[37499] = 16'hf72d;
  rom[37500] = 16'h62e4;
  rom[37501] = 16'hb573;
  rom[37502] = 16'hffff;
  rom[37503] = 16'hffff;
  rom[37504] = 16'hffff;
  rom[37505] = 16'hffff;
  rom[37506] = 16'hffff;
  rom[37507] = 16'hffff;
  rom[37508] = 16'hffff;
  rom[37509] = 16'hffff;
  rom[37510] = 16'hffff;
  rom[37511] = 16'hffff;
  rom[37512] = 16'hffff;
  rom[37513] = 16'hffff;
  rom[37514] = 16'hffff;
  rom[37515] = 16'hffff;
  rom[37516] = 16'hffff;
  rom[37517] = 16'hffff;
  rom[37518] = 16'hffff;
  rom[37519] = 16'hffff;
  rom[37520] = 16'hffff;
  rom[37521] = 16'hffff;
  rom[37522] = 16'hffff;
  rom[37523] = 16'hffff;
  rom[37524] = 16'hffff;
  rom[37525] = 16'hffff;
  rom[37526] = 16'hffff;
  rom[37527] = 16'hffff;
  rom[37528] = 16'hffff;
  rom[37529] = 16'hffff;
  rom[37530] = 16'hffff;
  rom[37531] = 16'hffff;
  rom[37532] = 16'hffff;
  rom[37533] = 16'hffff;
  rom[37534] = 16'hffff;
  rom[37535] = 16'hffff;
  rom[37536] = 16'hffff;
  rom[37537] = 16'hffff;
  rom[37538] = 16'hffff;
  rom[37539] = 16'hffff;
  rom[37540] = 16'hffff;
  rom[37541] = 16'hffff;
  rom[37542] = 16'hffff;
  rom[37543] = 16'hffff;
  rom[37544] = 16'hffff;
  rom[37545] = 16'hffff;
  rom[37546] = 16'hffff;
  rom[37547] = 16'hffff;
  rom[37548] = 16'hffff;
  rom[37549] = 16'hffff;
  rom[37550] = 16'hffff;
  rom[37551] = 16'hffff;
  rom[37552] = 16'hffff;
  rom[37553] = 16'hffff;
  rom[37554] = 16'hffff;
  rom[37555] = 16'hffff;
  rom[37556] = 16'hffff;
  rom[37557] = 16'hffff;
  rom[37558] = 16'hffff;
  rom[37559] = 16'hffff;
  rom[37560] = 16'hffff;
  rom[37561] = 16'hffff;
  rom[37562] = 16'hffff;
  rom[37563] = 16'hffff;
  rom[37564] = 16'hffff;
  rom[37565] = 16'hffff;
  rom[37566] = 16'hffff;
  rom[37567] = 16'hffff;
  rom[37568] = 16'hffff;
  rom[37569] = 16'hffff;
  rom[37570] = 16'hffff;
  rom[37571] = 16'hffff;
  rom[37572] = 16'hffff;
  rom[37573] = 16'hffff;
  rom[37574] = 16'hffff;
  rom[37575] = 16'hffff;
  rom[37576] = 16'hffff;
  rom[37577] = 16'hffff;
  rom[37578] = 16'hffff;
  rom[37579] = 16'hffff;
  rom[37580] = 16'hffff;
  rom[37581] = 16'hffff;
  rom[37582] = 16'hffff;
  rom[37583] = 16'hffff;
  rom[37584] = 16'hffff;
  rom[37585] = 16'hffff;
  rom[37586] = 16'hffff;
  rom[37587] = 16'hffff;
  rom[37588] = 16'hffff;
  rom[37589] = 16'hffff;
  rom[37590] = 16'hffff;
  rom[37591] = 16'hffff;
  rom[37592] = 16'hffff;
  rom[37593] = 16'hffff;
  rom[37594] = 16'hffff;
  rom[37595] = 16'hffff;
  rom[37596] = 16'hffff;
  rom[37597] = 16'hffff;
  rom[37598] = 16'hffff;
  rom[37599] = 16'hffff;
  rom[37600] = 16'hffff;
  rom[37601] = 16'hffff;
  rom[37602] = 16'hffff;
  rom[37603] = 16'hffff;
  rom[37604] = 16'hffff;
  rom[37605] = 16'hffff;
  rom[37606] = 16'hffff;
  rom[37607] = 16'hffff;
  rom[37608] = 16'hffff;
  rom[37609] = 16'hffff;
  rom[37610] = 16'hffff;
  rom[37611] = 16'hffff;
  rom[37612] = 16'hffff;
  rom[37613] = 16'hffff;
  rom[37614] = 16'hffff;
  rom[37615] = 16'hffff;
  rom[37616] = 16'hffff;
  rom[37617] = 16'hffff;
  rom[37618] = 16'hffff;
  rom[37619] = 16'hffff;
  rom[37620] = 16'hffff;
  rom[37621] = 16'hffff;
  rom[37622] = 16'hffff;
  rom[37623] = 16'hffff;
  rom[37624] = 16'hffff;
  rom[37625] = 16'hffff;
  rom[37626] = 16'hffff;
  rom[37627] = 16'hffff;
  rom[37628] = 16'hffff;
  rom[37629] = 16'hffff;
  rom[37630] = 16'hffff;
  rom[37631] = 16'hffff;
  rom[37632] = 16'hffff;
  rom[37633] = 16'hffff;
  rom[37634] = 16'hffff;
  rom[37635] = 16'hffff;
  rom[37636] = 16'hffff;
  rom[37637] = 16'hffff;
  rom[37638] = 16'hffff;
  rom[37639] = 16'hffff;
  rom[37640] = 16'hffff;
  rom[37641] = 16'hffff;
  rom[37642] = 16'hffff;
  rom[37643] = 16'hffff;
  rom[37644] = 16'hffff;
  rom[37645] = 16'hffff;
  rom[37646] = 16'hffff;
  rom[37647] = 16'hffff;
  rom[37648] = 16'hffff;
  rom[37649] = 16'hffff;
  rom[37650] = 16'hffff;
  rom[37651] = 16'hffff;
  rom[37652] = 16'hffff;
  rom[37653] = 16'hffff;
  rom[37654] = 16'hffff;
  rom[37655] = 16'hffff;
  rom[37656] = 16'hffff;
  rom[37657] = 16'hffff;
  rom[37658] = 16'hffff;
  rom[37659] = 16'hffff;
  rom[37660] = 16'hffff;
  rom[37661] = 16'hffff;
  rom[37662] = 16'hffff;
  rom[37663] = 16'hffff;
  rom[37664] = 16'hffff;
  rom[37665] = 16'hffff;
  rom[37666] = 16'hffff;
  rom[37667] = 16'hffff;
  rom[37668] = 16'hffff;
  rom[37669] = 16'hffff;
  rom[37670] = 16'hffff;
  rom[37671] = 16'hffff;
  rom[37672] = 16'hffff;
  rom[37673] = 16'hffff;
  rom[37674] = 16'hffff;
  rom[37675] = 16'hffff;
  rom[37676] = 16'hffdd;
  rom[37677] = 16'h7368;
  rom[37678] = 16'hb58b;
  rom[37679] = 16'hf72d;
  rom[37680] = 16'hf70a;
  rom[37681] = 16'hff49;
  rom[37682] = 16'hf727;
  rom[37683] = 16'hff48;
  rom[37684] = 16'hf708;
  rom[37685] = 16'hff28;
  rom[37686] = 16'hff08;
  rom[37687] = 16'hff28;
  rom[37688] = 16'hf708;
  rom[37689] = 16'hff28;
  rom[37690] = 16'hff08;
  rom[37691] = 16'hff29;
  rom[37692] = 16'hf709;
  rom[37693] = 16'hf729;
  rom[37694] = 16'hf708;
  rom[37695] = 16'hff28;
  rom[37696] = 16'hf708;
  rom[37697] = 16'hff2a;
  rom[37698] = 16'hff2a;
  rom[37699] = 16'he68b;
  rom[37700] = 16'h4a21;
  rom[37701] = 16'hd677;
  rom[37702] = 16'hffde;
  rom[37703] = 16'hffff;
  rom[37704] = 16'hffff;
  rom[37705] = 16'hffff;
  rom[37706] = 16'hffff;
  rom[37707] = 16'hffff;
  rom[37708] = 16'hffff;
  rom[37709] = 16'hffff;
  rom[37710] = 16'hffff;
  rom[37711] = 16'hffff;
  rom[37712] = 16'hffff;
  rom[37713] = 16'hffff;
  rom[37714] = 16'hffff;
  rom[37715] = 16'hffff;
  rom[37716] = 16'hffff;
  rom[37717] = 16'hffff;
  rom[37718] = 16'hffff;
  rom[37719] = 16'hffff;
  rom[37720] = 16'hffff;
  rom[37721] = 16'hffff;
  rom[37722] = 16'hffff;
  rom[37723] = 16'hffff;
  rom[37724] = 16'hffff;
  rom[37725] = 16'hffff;
  rom[37726] = 16'hffff;
  rom[37727] = 16'hffff;
  rom[37728] = 16'hffff;
  rom[37729] = 16'hffff;
  rom[37730] = 16'hffff;
  rom[37731] = 16'hffff;
  rom[37732] = 16'hffff;
  rom[37733] = 16'hffff;
  rom[37734] = 16'hffff;
  rom[37735] = 16'hffff;
  rom[37736] = 16'hffff;
  rom[37737] = 16'hffff;
  rom[37738] = 16'hffff;
  rom[37739] = 16'hffff;
  rom[37740] = 16'hffff;
  rom[37741] = 16'hffff;
  rom[37742] = 16'hffff;
  rom[37743] = 16'hffff;
  rom[37744] = 16'hffff;
  rom[37745] = 16'hffff;
  rom[37746] = 16'hffff;
  rom[37747] = 16'hffff;
  rom[37748] = 16'hffff;
  rom[37749] = 16'hffff;
  rom[37750] = 16'hffff;
  rom[37751] = 16'hffff;
  rom[37752] = 16'hffff;
  rom[37753] = 16'hffff;
  rom[37754] = 16'hffff;
  rom[37755] = 16'hffff;
  rom[37756] = 16'hffff;
  rom[37757] = 16'hffff;
  rom[37758] = 16'hffff;
  rom[37759] = 16'hffff;
  rom[37760] = 16'hffff;
  rom[37761] = 16'hffff;
  rom[37762] = 16'hffff;
  rom[37763] = 16'hffff;
  rom[37764] = 16'hffff;
  rom[37765] = 16'hffff;
  rom[37766] = 16'hffff;
  rom[37767] = 16'hffff;
  rom[37768] = 16'hffff;
  rom[37769] = 16'hffff;
  rom[37770] = 16'hffff;
  rom[37771] = 16'hffff;
  rom[37772] = 16'hffff;
  rom[37773] = 16'hffff;
  rom[37774] = 16'hffff;
  rom[37775] = 16'hffff;
  rom[37776] = 16'hffff;
  rom[37777] = 16'hffff;
  rom[37778] = 16'hffff;
  rom[37779] = 16'hffff;
  rom[37780] = 16'hffff;
  rom[37781] = 16'hffff;
  rom[37782] = 16'hffff;
  rom[37783] = 16'hffff;
  rom[37784] = 16'hffff;
  rom[37785] = 16'hffff;
  rom[37786] = 16'hffff;
  rom[37787] = 16'hffff;
  rom[37788] = 16'hffff;
  rom[37789] = 16'hffff;
  rom[37790] = 16'hffff;
  rom[37791] = 16'hffff;
  rom[37792] = 16'hffff;
  rom[37793] = 16'hffff;
  rom[37794] = 16'hffff;
  rom[37795] = 16'hffff;
  rom[37796] = 16'hffff;
  rom[37797] = 16'hffff;
  rom[37798] = 16'hffff;
  rom[37799] = 16'hffff;
  rom[37800] = 16'hffff;
  rom[37801] = 16'hffff;
  rom[37802] = 16'hffff;
  rom[37803] = 16'hffff;
  rom[37804] = 16'hffff;
  rom[37805] = 16'hffff;
  rom[37806] = 16'hffff;
  rom[37807] = 16'hffff;
  rom[37808] = 16'hffff;
  rom[37809] = 16'hffff;
  rom[37810] = 16'hffff;
  rom[37811] = 16'hffff;
  rom[37812] = 16'hffff;
  rom[37813] = 16'hffff;
  rom[37814] = 16'hffff;
  rom[37815] = 16'hffff;
  rom[37816] = 16'hffff;
  rom[37817] = 16'hffff;
  rom[37818] = 16'hffff;
  rom[37819] = 16'hffff;
  rom[37820] = 16'hffff;
  rom[37821] = 16'hffff;
  rom[37822] = 16'hffff;
  rom[37823] = 16'hffff;
  rom[37824] = 16'hffff;
  rom[37825] = 16'hffff;
  rom[37826] = 16'hffff;
  rom[37827] = 16'hffff;
  rom[37828] = 16'hffff;
  rom[37829] = 16'hffff;
  rom[37830] = 16'hffff;
  rom[37831] = 16'hffff;
  rom[37832] = 16'hffff;
  rom[37833] = 16'hffff;
  rom[37834] = 16'hffff;
  rom[37835] = 16'hffff;
  rom[37836] = 16'hffff;
  rom[37837] = 16'hffff;
  rom[37838] = 16'hffff;
  rom[37839] = 16'hffff;
  rom[37840] = 16'hffff;
  rom[37841] = 16'hffff;
  rom[37842] = 16'hffff;
  rom[37843] = 16'hffff;
  rom[37844] = 16'hffff;
  rom[37845] = 16'hffff;
  rom[37846] = 16'hffff;
  rom[37847] = 16'hffff;
  rom[37848] = 16'hffff;
  rom[37849] = 16'hffff;
  rom[37850] = 16'hffff;
  rom[37851] = 16'hffff;
  rom[37852] = 16'hffff;
  rom[37853] = 16'hffff;
  rom[37854] = 16'hffff;
  rom[37855] = 16'hffff;
  rom[37856] = 16'hffff;
  rom[37857] = 16'hffff;
  rom[37858] = 16'hffff;
  rom[37859] = 16'hffff;
  rom[37860] = 16'hffff;
  rom[37861] = 16'hffff;
  rom[37862] = 16'hffff;
  rom[37863] = 16'hffff;
  rom[37864] = 16'hffff;
  rom[37865] = 16'hffff;
  rom[37866] = 16'hffff;
  rom[37867] = 16'hffff;
  rom[37868] = 16'hffff;
  rom[37869] = 16'hffff;
  rom[37870] = 16'hffff;
  rom[37871] = 16'hffff;
  rom[37872] = 16'hffff;
  rom[37873] = 16'hffff;
  rom[37874] = 16'hffff;
  rom[37875] = 16'hffff;
  rom[37876] = 16'hfffe;
  rom[37877] = 16'hb572;
  rom[37878] = 16'h7345;
  rom[37879] = 16'heeee;
  rom[37880] = 16'hf70b;
  rom[37881] = 16'hf74a;
  rom[37882] = 16'hff48;
  rom[37883] = 16'hf728;
  rom[37884] = 16'hff49;
  rom[37885] = 16'hff28;
  rom[37886] = 16'hff29;
  rom[37887] = 16'hff28;
  rom[37888] = 16'hff29;
  rom[37889] = 16'hff29;
  rom[37890] = 16'hff29;
  rom[37891] = 16'hff28;
  rom[37892] = 16'hff2a;
  rom[37893] = 16'hf729;
  rom[37894] = 16'hff29;
  rom[37895] = 16'hff28;
  rom[37896] = 16'hff2a;
  rom[37897] = 16'hff09;
  rom[37898] = 16'hff0a;
  rom[37899] = 16'hde6a;
  rom[37900] = 16'h5a62;
  rom[37901] = 16'hde98;
  rom[37902] = 16'hffff;
  rom[37903] = 16'hffff;
  rom[37904] = 16'hffff;
  rom[37905] = 16'hffff;
  rom[37906] = 16'hffff;
  rom[37907] = 16'hffff;
  rom[37908] = 16'hffff;
  rom[37909] = 16'hffff;
  rom[37910] = 16'hffff;
  rom[37911] = 16'hffff;
  rom[37912] = 16'hffff;
  rom[37913] = 16'hffff;
  rom[37914] = 16'hffff;
  rom[37915] = 16'hffff;
  rom[37916] = 16'hffff;
  rom[37917] = 16'hffff;
  rom[37918] = 16'hffff;
  rom[37919] = 16'hffff;
  rom[37920] = 16'hffff;
  rom[37921] = 16'hffff;
  rom[37922] = 16'hffff;
  rom[37923] = 16'hffff;
  rom[37924] = 16'hffff;
  rom[37925] = 16'hffff;
  rom[37926] = 16'hffff;
  rom[37927] = 16'hffff;
  rom[37928] = 16'hffff;
  rom[37929] = 16'hffff;
  rom[37930] = 16'hffff;
  rom[37931] = 16'hffff;
  rom[37932] = 16'hffff;
  rom[37933] = 16'hffff;
  rom[37934] = 16'hffff;
  rom[37935] = 16'hffff;
  rom[37936] = 16'hffff;
  rom[37937] = 16'hffff;
  rom[37938] = 16'hffff;
  rom[37939] = 16'hffff;
  rom[37940] = 16'hffff;
  rom[37941] = 16'hffff;
  rom[37942] = 16'hffff;
  rom[37943] = 16'hffff;
  rom[37944] = 16'hffff;
  rom[37945] = 16'hffff;
  rom[37946] = 16'hffff;
  rom[37947] = 16'hffff;
  rom[37948] = 16'hffff;
  rom[37949] = 16'hffff;
  rom[37950] = 16'hffff;
  rom[37951] = 16'hffff;
  rom[37952] = 16'hffff;
  rom[37953] = 16'hffff;
  rom[37954] = 16'hffff;
  rom[37955] = 16'hffff;
  rom[37956] = 16'hffff;
  rom[37957] = 16'hffff;
  rom[37958] = 16'hffff;
  rom[37959] = 16'hffff;
  rom[37960] = 16'hffff;
  rom[37961] = 16'hffff;
  rom[37962] = 16'hffff;
  rom[37963] = 16'hffff;
  rom[37964] = 16'hffff;
  rom[37965] = 16'hffff;
  rom[37966] = 16'hffff;
  rom[37967] = 16'hffff;
  rom[37968] = 16'hffff;
  rom[37969] = 16'hffff;
  rom[37970] = 16'hffff;
  rom[37971] = 16'hffff;
  rom[37972] = 16'hffff;
  rom[37973] = 16'hffff;
  rom[37974] = 16'hffff;
  rom[37975] = 16'hffff;
  rom[37976] = 16'hffff;
  rom[37977] = 16'hffff;
  rom[37978] = 16'hffff;
  rom[37979] = 16'hffff;
  rom[37980] = 16'hffff;
  rom[37981] = 16'hffff;
  rom[37982] = 16'hffff;
  rom[37983] = 16'hffff;
  rom[37984] = 16'hffff;
  rom[37985] = 16'hffff;
  rom[37986] = 16'hffff;
  rom[37987] = 16'hffff;
  rom[37988] = 16'hffff;
  rom[37989] = 16'hffff;
  rom[37990] = 16'hffff;
  rom[37991] = 16'hffff;
  rom[37992] = 16'hffff;
  rom[37993] = 16'hffff;
  rom[37994] = 16'hffff;
  rom[37995] = 16'hffff;
  rom[37996] = 16'hffff;
  rom[37997] = 16'hffff;
  rom[37998] = 16'hffff;
  rom[37999] = 16'hffff;
  rom[38000] = 16'hffff;
  rom[38001] = 16'hffff;
  rom[38002] = 16'hffff;
  rom[38003] = 16'hffff;
  rom[38004] = 16'hffff;
  rom[38005] = 16'hffff;
  rom[38006] = 16'hffff;
  rom[38007] = 16'hffff;
  rom[38008] = 16'hffff;
  rom[38009] = 16'hffff;
  rom[38010] = 16'hffff;
  rom[38011] = 16'hffff;
  rom[38012] = 16'hffff;
  rom[38013] = 16'hffff;
  rom[38014] = 16'hffff;
  rom[38015] = 16'hffff;
  rom[38016] = 16'hffff;
  rom[38017] = 16'hffff;
  rom[38018] = 16'hffff;
  rom[38019] = 16'hffff;
  rom[38020] = 16'hffff;
  rom[38021] = 16'hffff;
  rom[38022] = 16'hffff;
  rom[38023] = 16'hffff;
  rom[38024] = 16'hffff;
  rom[38025] = 16'hffff;
  rom[38026] = 16'hffff;
  rom[38027] = 16'hffff;
  rom[38028] = 16'hffff;
  rom[38029] = 16'hffff;
  rom[38030] = 16'hffff;
  rom[38031] = 16'hffff;
  rom[38032] = 16'hffff;
  rom[38033] = 16'hffff;
  rom[38034] = 16'hffff;
  rom[38035] = 16'hffff;
  rom[38036] = 16'hffff;
  rom[38037] = 16'hffff;
  rom[38038] = 16'hffff;
  rom[38039] = 16'hffff;
  rom[38040] = 16'hffff;
  rom[38041] = 16'hffff;
  rom[38042] = 16'hffff;
  rom[38043] = 16'hffff;
  rom[38044] = 16'hffff;
  rom[38045] = 16'hffff;
  rom[38046] = 16'hffff;
  rom[38047] = 16'hffff;
  rom[38048] = 16'hffff;
  rom[38049] = 16'hffff;
  rom[38050] = 16'hffff;
  rom[38051] = 16'hffff;
  rom[38052] = 16'hffff;
  rom[38053] = 16'hffff;
  rom[38054] = 16'hffff;
  rom[38055] = 16'hffff;
  rom[38056] = 16'hffff;
  rom[38057] = 16'hffff;
  rom[38058] = 16'hffff;
  rom[38059] = 16'hffff;
  rom[38060] = 16'hffff;
  rom[38061] = 16'hffff;
  rom[38062] = 16'hffff;
  rom[38063] = 16'hffff;
  rom[38064] = 16'hffff;
  rom[38065] = 16'hffff;
  rom[38066] = 16'hffff;
  rom[38067] = 16'hffff;
  rom[38068] = 16'hffff;
  rom[38069] = 16'hffff;
  rom[38070] = 16'hffff;
  rom[38071] = 16'hffff;
  rom[38072] = 16'hffff;
  rom[38073] = 16'hffff;
  rom[38074] = 16'hffff;
  rom[38075] = 16'hffff;
  rom[38076] = 16'hffde;
  rom[38077] = 16'hdeb9;
  rom[38078] = 16'h4a03;
  rom[38079] = 16'heeef;
  rom[38080] = 16'hf72c;
  rom[38081] = 16'hf709;
  rom[38082] = 16'hf728;
  rom[38083] = 16'hf728;
  rom[38084] = 16'hff28;
  rom[38085] = 16'hff29;
  rom[38086] = 16'hf709;
  rom[38087] = 16'hff29;
  rom[38088] = 16'hff09;
  rom[38089] = 16'hff29;
  rom[38090] = 16'hf708;
  rom[38091] = 16'hff29;
  rom[38092] = 16'hf709;
  rom[38093] = 16'hf729;
  rom[38094] = 16'hf728;
  rom[38095] = 16'hff28;
  rom[38096] = 16'hfee9;
  rom[38097] = 16'hfee9;
  rom[38098] = 16'hf6ea;
  rom[38099] = 16'hd62a;
  rom[38100] = 16'h5242;
  rom[38101] = 16'hdeb8;
  rom[38102] = 16'hffff;
  rom[38103] = 16'hffff;
  rom[38104] = 16'hffff;
  rom[38105] = 16'hffff;
  rom[38106] = 16'hffff;
  rom[38107] = 16'hffff;
  rom[38108] = 16'hffff;
  rom[38109] = 16'hffff;
  rom[38110] = 16'hffff;
  rom[38111] = 16'hffff;
  rom[38112] = 16'hffff;
  rom[38113] = 16'hffff;
  rom[38114] = 16'hffff;
  rom[38115] = 16'hffff;
  rom[38116] = 16'hffff;
  rom[38117] = 16'hffff;
  rom[38118] = 16'hffff;
  rom[38119] = 16'hffff;
  rom[38120] = 16'hffff;
  rom[38121] = 16'hffff;
  rom[38122] = 16'hffff;
  rom[38123] = 16'hffff;
  rom[38124] = 16'hffff;
  rom[38125] = 16'hffff;
  rom[38126] = 16'hffff;
  rom[38127] = 16'hffff;
  rom[38128] = 16'hffff;
  rom[38129] = 16'hffff;
  rom[38130] = 16'hffff;
  rom[38131] = 16'hffff;
  rom[38132] = 16'hffff;
  rom[38133] = 16'hffff;
  rom[38134] = 16'hffff;
  rom[38135] = 16'hffff;
  rom[38136] = 16'hffff;
  rom[38137] = 16'hffff;
  rom[38138] = 16'hffff;
  rom[38139] = 16'hffff;
  rom[38140] = 16'hffff;
  rom[38141] = 16'hffff;
  rom[38142] = 16'hffff;
  rom[38143] = 16'hffff;
  rom[38144] = 16'hffff;
  rom[38145] = 16'hffff;
  rom[38146] = 16'hffff;
  rom[38147] = 16'hffff;
  rom[38148] = 16'hffff;
  rom[38149] = 16'hffff;
  rom[38150] = 16'hffff;
  rom[38151] = 16'hffff;
  rom[38152] = 16'hffff;
  rom[38153] = 16'hffff;
  rom[38154] = 16'hffff;
  rom[38155] = 16'hffff;
  rom[38156] = 16'hffff;
  rom[38157] = 16'hffff;
  rom[38158] = 16'hffff;
  rom[38159] = 16'hffff;
  rom[38160] = 16'hffff;
  rom[38161] = 16'hffff;
  rom[38162] = 16'hffff;
  rom[38163] = 16'hffff;
  rom[38164] = 16'hffff;
  rom[38165] = 16'hffff;
  rom[38166] = 16'hffff;
  rom[38167] = 16'hffff;
  rom[38168] = 16'hffff;
  rom[38169] = 16'hffff;
  rom[38170] = 16'hffff;
  rom[38171] = 16'hffff;
  rom[38172] = 16'hffff;
  rom[38173] = 16'hffff;
  rom[38174] = 16'hffff;
  rom[38175] = 16'hffff;
  rom[38176] = 16'hffff;
  rom[38177] = 16'hffff;
  rom[38178] = 16'hffff;
  rom[38179] = 16'hffff;
  rom[38180] = 16'hffff;
  rom[38181] = 16'hffff;
  rom[38182] = 16'hffff;
  rom[38183] = 16'hffff;
  rom[38184] = 16'hffff;
  rom[38185] = 16'hffff;
  rom[38186] = 16'hffff;
  rom[38187] = 16'hffff;
  rom[38188] = 16'hffff;
  rom[38189] = 16'hffff;
  rom[38190] = 16'hffff;
  rom[38191] = 16'hffff;
  rom[38192] = 16'hffff;
  rom[38193] = 16'hffff;
  rom[38194] = 16'hffff;
  rom[38195] = 16'hffff;
  rom[38196] = 16'hffff;
  rom[38197] = 16'hffff;
  rom[38198] = 16'hffff;
  rom[38199] = 16'hffff;
  rom[38200] = 16'hffff;
  rom[38201] = 16'hffff;
  rom[38202] = 16'hffff;
  rom[38203] = 16'hffff;
  rom[38204] = 16'hffff;
  rom[38205] = 16'hffff;
  rom[38206] = 16'hffff;
  rom[38207] = 16'hffff;
  rom[38208] = 16'hffff;
  rom[38209] = 16'hffff;
  rom[38210] = 16'hffff;
  rom[38211] = 16'hffff;
  rom[38212] = 16'hffff;
  rom[38213] = 16'hffff;
  rom[38214] = 16'hffff;
  rom[38215] = 16'hffff;
  rom[38216] = 16'hffff;
  rom[38217] = 16'hffff;
  rom[38218] = 16'hffff;
  rom[38219] = 16'hffff;
  rom[38220] = 16'hffff;
  rom[38221] = 16'hffff;
  rom[38222] = 16'hffff;
  rom[38223] = 16'hffff;
  rom[38224] = 16'hffff;
  rom[38225] = 16'hffff;
  rom[38226] = 16'hffff;
  rom[38227] = 16'hffff;
  rom[38228] = 16'hffff;
  rom[38229] = 16'hffff;
  rom[38230] = 16'hffff;
  rom[38231] = 16'hffff;
  rom[38232] = 16'hffff;
  rom[38233] = 16'hffff;
  rom[38234] = 16'hffff;
  rom[38235] = 16'hffff;
  rom[38236] = 16'hffff;
  rom[38237] = 16'hffff;
  rom[38238] = 16'hffff;
  rom[38239] = 16'hffff;
  rom[38240] = 16'hffff;
  rom[38241] = 16'hffff;
  rom[38242] = 16'hffff;
  rom[38243] = 16'hffff;
  rom[38244] = 16'hffff;
  rom[38245] = 16'hffff;
  rom[38246] = 16'hffff;
  rom[38247] = 16'hffff;
  rom[38248] = 16'hffff;
  rom[38249] = 16'hffff;
  rom[38250] = 16'hffff;
  rom[38251] = 16'hffff;
  rom[38252] = 16'hffff;
  rom[38253] = 16'hffff;
  rom[38254] = 16'hffff;
  rom[38255] = 16'hffff;
  rom[38256] = 16'hffff;
  rom[38257] = 16'hffff;
  rom[38258] = 16'hffff;
  rom[38259] = 16'hffff;
  rom[38260] = 16'hffff;
  rom[38261] = 16'hffff;
  rom[38262] = 16'hffff;
  rom[38263] = 16'hffff;
  rom[38264] = 16'hffff;
  rom[38265] = 16'hffff;
  rom[38266] = 16'hffff;
  rom[38267] = 16'hffff;
  rom[38268] = 16'hffff;
  rom[38269] = 16'hffff;
  rom[38270] = 16'hffff;
  rom[38271] = 16'hffff;
  rom[38272] = 16'hffff;
  rom[38273] = 16'hffff;
  rom[38274] = 16'hffff;
  rom[38275] = 16'hffff;
  rom[38276] = 16'hffff;
  rom[38277] = 16'hffbe;
  rom[38278] = 16'h6b09;
  rom[38279] = 16'h9426;
  rom[38280] = 16'hf6ec;
  rom[38281] = 16'hff2a;
  rom[38282] = 16'hff29;
  rom[38283] = 16'hff4a;
  rom[38284] = 16'hff09;
  rom[38285] = 16'hff29;
  rom[38286] = 16'hff29;
  rom[38287] = 16'hff29;
  rom[38288] = 16'hff2a;
  rom[38289] = 16'hff09;
  rom[38290] = 16'hff29;
  rom[38291] = 16'hff28;
  rom[38292] = 16'hff29;
  rom[38293] = 16'hf729;
  rom[38294] = 16'hff29;
  rom[38295] = 16'hff28;
  rom[38296] = 16'hff0a;
  rom[38297] = 16'hfee9;
  rom[38298] = 16'hff2b;
  rom[38299] = 16'hcde9;
  rom[38300] = 16'h5242;
  rom[38301] = 16'he6d9;
  rom[38302] = 16'hffff;
  rom[38303] = 16'hffff;
  rom[38304] = 16'hffff;
  rom[38305] = 16'hffff;
  rom[38306] = 16'hffff;
  rom[38307] = 16'hffff;
  rom[38308] = 16'hffff;
  rom[38309] = 16'hffff;
  rom[38310] = 16'hffff;
  rom[38311] = 16'hffff;
  rom[38312] = 16'hffff;
  rom[38313] = 16'hffff;
  rom[38314] = 16'hffff;
  rom[38315] = 16'hffff;
  rom[38316] = 16'hffff;
  rom[38317] = 16'hffff;
  rom[38318] = 16'hffff;
  rom[38319] = 16'hffff;
  rom[38320] = 16'hffff;
  rom[38321] = 16'hffff;
  rom[38322] = 16'hffff;
  rom[38323] = 16'hffff;
  rom[38324] = 16'hffff;
  rom[38325] = 16'hffff;
  rom[38326] = 16'hffff;
  rom[38327] = 16'hffff;
  rom[38328] = 16'hffff;
  rom[38329] = 16'hffff;
  rom[38330] = 16'hffff;
  rom[38331] = 16'hffff;
  rom[38332] = 16'hffff;
  rom[38333] = 16'hffff;
  rom[38334] = 16'hffff;
  rom[38335] = 16'hffff;
  rom[38336] = 16'hffff;
  rom[38337] = 16'hffff;
  rom[38338] = 16'hffff;
  rom[38339] = 16'hffff;
  rom[38340] = 16'hffff;
  rom[38341] = 16'hffff;
  rom[38342] = 16'hffff;
  rom[38343] = 16'hffff;
  rom[38344] = 16'hffff;
  rom[38345] = 16'hffff;
  rom[38346] = 16'hffff;
  rom[38347] = 16'hffff;
  rom[38348] = 16'hffff;
  rom[38349] = 16'hffff;
  rom[38350] = 16'hffff;
  rom[38351] = 16'hffff;
  rom[38352] = 16'hffff;
  rom[38353] = 16'hffff;
  rom[38354] = 16'hffff;
  rom[38355] = 16'hffff;
  rom[38356] = 16'hffff;
  rom[38357] = 16'hffff;
  rom[38358] = 16'hffff;
  rom[38359] = 16'hffff;
  rom[38360] = 16'hffff;
  rom[38361] = 16'hffff;
  rom[38362] = 16'hffff;
  rom[38363] = 16'hffff;
  rom[38364] = 16'hffff;
  rom[38365] = 16'hffff;
  rom[38366] = 16'hffff;
  rom[38367] = 16'hffff;
  rom[38368] = 16'hffff;
  rom[38369] = 16'hffff;
  rom[38370] = 16'hffff;
  rom[38371] = 16'hffff;
  rom[38372] = 16'hffff;
  rom[38373] = 16'hffff;
  rom[38374] = 16'hffff;
  rom[38375] = 16'hffff;
  rom[38376] = 16'hffff;
  rom[38377] = 16'hffff;
  rom[38378] = 16'hffff;
  rom[38379] = 16'hffff;
  rom[38380] = 16'hffff;
  rom[38381] = 16'hffff;
  rom[38382] = 16'hffff;
  rom[38383] = 16'hffff;
  rom[38384] = 16'hffff;
  rom[38385] = 16'hffff;
  rom[38386] = 16'hffff;
  rom[38387] = 16'hffff;
  rom[38388] = 16'hffff;
  rom[38389] = 16'hffff;
  rom[38390] = 16'hffff;
  rom[38391] = 16'hffff;
  rom[38392] = 16'hffff;
  rom[38393] = 16'hffff;
  rom[38394] = 16'hffff;
  rom[38395] = 16'hffff;
  rom[38396] = 16'hffff;
  rom[38397] = 16'hffff;
  rom[38398] = 16'hffff;
  rom[38399] = 16'hffff;
  rom[38400] = 16'hffff;
  rom[38401] = 16'hffff;
  rom[38402] = 16'hffff;
  rom[38403] = 16'hffff;
  rom[38404] = 16'hffff;
  rom[38405] = 16'hffff;
  rom[38406] = 16'hffff;
  rom[38407] = 16'hffff;
  rom[38408] = 16'hffff;
  rom[38409] = 16'hffff;
  rom[38410] = 16'hffff;
  rom[38411] = 16'hffff;
  rom[38412] = 16'hffff;
  rom[38413] = 16'hffff;
  rom[38414] = 16'hffff;
  rom[38415] = 16'hffff;
  rom[38416] = 16'hffff;
  rom[38417] = 16'hffff;
  rom[38418] = 16'hffff;
  rom[38419] = 16'hffff;
  rom[38420] = 16'hffff;
  rom[38421] = 16'hffff;
  rom[38422] = 16'hffff;
  rom[38423] = 16'hffff;
  rom[38424] = 16'hffff;
  rom[38425] = 16'hffff;
  rom[38426] = 16'hffff;
  rom[38427] = 16'hffff;
  rom[38428] = 16'hffff;
  rom[38429] = 16'hffff;
  rom[38430] = 16'hffff;
  rom[38431] = 16'hffff;
  rom[38432] = 16'hffff;
  rom[38433] = 16'hffff;
  rom[38434] = 16'hffff;
  rom[38435] = 16'hffff;
  rom[38436] = 16'hffff;
  rom[38437] = 16'hffff;
  rom[38438] = 16'hffff;
  rom[38439] = 16'hffff;
  rom[38440] = 16'hffff;
  rom[38441] = 16'hffff;
  rom[38442] = 16'hffff;
  rom[38443] = 16'hffff;
  rom[38444] = 16'hffff;
  rom[38445] = 16'hffff;
  rom[38446] = 16'hffff;
  rom[38447] = 16'hffff;
  rom[38448] = 16'hffff;
  rom[38449] = 16'hffff;
  rom[38450] = 16'hffff;
  rom[38451] = 16'hffff;
  rom[38452] = 16'hffff;
  rom[38453] = 16'hffff;
  rom[38454] = 16'hffff;
  rom[38455] = 16'hffff;
  rom[38456] = 16'hffff;
  rom[38457] = 16'hffff;
  rom[38458] = 16'hffff;
  rom[38459] = 16'hffff;
  rom[38460] = 16'hffff;
  rom[38461] = 16'hffff;
  rom[38462] = 16'hffff;
  rom[38463] = 16'hffff;
  rom[38464] = 16'hffff;
  rom[38465] = 16'hffff;
  rom[38466] = 16'hffff;
  rom[38467] = 16'hffff;
  rom[38468] = 16'hffff;
  rom[38469] = 16'hffff;
  rom[38470] = 16'hffff;
  rom[38471] = 16'hffff;
  rom[38472] = 16'hffff;
  rom[38473] = 16'hffff;
  rom[38474] = 16'hffff;
  rom[38475] = 16'hffff;
  rom[38476] = 16'hffde;
  rom[38477] = 16'hffff;
  rom[38478] = 16'hb553;
  rom[38479] = 16'h5a82;
  rom[38480] = 16'hde8b;
  rom[38481] = 16'hff2a;
  rom[38482] = 16'hff09;
  rom[38483] = 16'hff0a;
  rom[38484] = 16'hf70a;
  rom[38485] = 16'hff29;
  rom[38486] = 16'hff28;
  rom[38487] = 16'hff09;
  rom[38488] = 16'hf709;
  rom[38489] = 16'hf729;
  rom[38490] = 16'hf728;
  rom[38491] = 16'hf748;
  rom[38492] = 16'hf728;
  rom[38493] = 16'hff29;
  rom[38494] = 16'hff08;
  rom[38495] = 16'hff29;
  rom[38496] = 16'hf709;
  rom[38497] = 16'hf709;
  rom[38498] = 16'hf70b;
  rom[38499] = 16'hcdaa;
  rom[38500] = 16'h4a01;
  rom[38501] = 16'he6fa;
  rom[38502] = 16'hffff;
  rom[38503] = 16'hffff;
  rom[38504] = 16'hffff;
  rom[38505] = 16'hffff;
  rom[38506] = 16'hffff;
  rom[38507] = 16'hffff;
  rom[38508] = 16'hffff;
  rom[38509] = 16'hffff;
  rom[38510] = 16'hffff;
  rom[38511] = 16'hffff;
  rom[38512] = 16'hffff;
  rom[38513] = 16'hffff;
  rom[38514] = 16'hffff;
  rom[38515] = 16'hffff;
  rom[38516] = 16'hffff;
  rom[38517] = 16'hffff;
  rom[38518] = 16'hffff;
  rom[38519] = 16'hffff;
  rom[38520] = 16'hffff;
  rom[38521] = 16'hffff;
  rom[38522] = 16'hffff;
  rom[38523] = 16'hffff;
  rom[38524] = 16'hffff;
  rom[38525] = 16'hffff;
  rom[38526] = 16'hffff;
  rom[38527] = 16'hffff;
  rom[38528] = 16'hffff;
  rom[38529] = 16'hffff;
  rom[38530] = 16'hffff;
  rom[38531] = 16'hffff;
  rom[38532] = 16'hffff;
  rom[38533] = 16'hffff;
  rom[38534] = 16'hffff;
  rom[38535] = 16'hffff;
  rom[38536] = 16'hffff;
  rom[38537] = 16'hffff;
  rom[38538] = 16'hffff;
  rom[38539] = 16'hffff;
  rom[38540] = 16'hffff;
  rom[38541] = 16'hffff;
  rom[38542] = 16'hffff;
  rom[38543] = 16'hffff;
  rom[38544] = 16'hffff;
  rom[38545] = 16'hffff;
  rom[38546] = 16'hffff;
  rom[38547] = 16'hffff;
  rom[38548] = 16'hffff;
  rom[38549] = 16'hffff;
  rom[38550] = 16'hffff;
  rom[38551] = 16'hffff;
  rom[38552] = 16'hffff;
  rom[38553] = 16'hffff;
  rom[38554] = 16'hffff;
  rom[38555] = 16'hffff;
  rom[38556] = 16'hffff;
  rom[38557] = 16'hffff;
  rom[38558] = 16'hffff;
  rom[38559] = 16'hffff;
  rom[38560] = 16'hffff;
  rom[38561] = 16'hffff;
  rom[38562] = 16'hffff;
  rom[38563] = 16'hffff;
  rom[38564] = 16'hffff;
  rom[38565] = 16'hffff;
  rom[38566] = 16'hffff;
  rom[38567] = 16'hffff;
  rom[38568] = 16'hffff;
  rom[38569] = 16'hffff;
  rom[38570] = 16'hffff;
  rom[38571] = 16'hffff;
  rom[38572] = 16'hffff;
  rom[38573] = 16'hffff;
  rom[38574] = 16'hffff;
  rom[38575] = 16'hffff;
  rom[38576] = 16'hffff;
  rom[38577] = 16'hffff;
  rom[38578] = 16'hffff;
  rom[38579] = 16'hffff;
  rom[38580] = 16'hffff;
  rom[38581] = 16'hffff;
  rom[38582] = 16'hffff;
  rom[38583] = 16'hffff;
  rom[38584] = 16'hffff;
  rom[38585] = 16'hffff;
  rom[38586] = 16'hffff;
  rom[38587] = 16'hffff;
  rom[38588] = 16'hffff;
  rom[38589] = 16'hffff;
  rom[38590] = 16'hffff;
  rom[38591] = 16'hffff;
  rom[38592] = 16'hffff;
  rom[38593] = 16'hffff;
  rom[38594] = 16'hffff;
  rom[38595] = 16'hffff;
  rom[38596] = 16'hffff;
  rom[38597] = 16'hffff;
  rom[38598] = 16'hffff;
  rom[38599] = 16'hffff;
  rom[38600] = 16'hffff;
  rom[38601] = 16'hffff;
  rom[38602] = 16'hffff;
  rom[38603] = 16'hffff;
  rom[38604] = 16'hffff;
  rom[38605] = 16'hffff;
  rom[38606] = 16'hffff;
  rom[38607] = 16'hffff;
  rom[38608] = 16'hffff;
  rom[38609] = 16'hffff;
  rom[38610] = 16'hffff;
  rom[38611] = 16'hffff;
  rom[38612] = 16'hffff;
  rom[38613] = 16'hffff;
  rom[38614] = 16'hffff;
  rom[38615] = 16'hffff;
  rom[38616] = 16'hffff;
  rom[38617] = 16'hffff;
  rom[38618] = 16'hffff;
  rom[38619] = 16'hffff;
  rom[38620] = 16'hffff;
  rom[38621] = 16'hffff;
  rom[38622] = 16'hffff;
  rom[38623] = 16'hffff;
  rom[38624] = 16'hffff;
  rom[38625] = 16'hffff;
  rom[38626] = 16'hffff;
  rom[38627] = 16'hffff;
  rom[38628] = 16'hffff;
  rom[38629] = 16'hffff;
  rom[38630] = 16'hffff;
  rom[38631] = 16'hffff;
  rom[38632] = 16'hffff;
  rom[38633] = 16'hffff;
  rom[38634] = 16'hffff;
  rom[38635] = 16'hffff;
  rom[38636] = 16'hffff;
  rom[38637] = 16'hffff;
  rom[38638] = 16'hffff;
  rom[38639] = 16'hffff;
  rom[38640] = 16'hffff;
  rom[38641] = 16'hffff;
  rom[38642] = 16'hffff;
  rom[38643] = 16'hffff;
  rom[38644] = 16'hffff;
  rom[38645] = 16'hffff;
  rom[38646] = 16'hffff;
  rom[38647] = 16'hffff;
  rom[38648] = 16'hffff;
  rom[38649] = 16'hffff;
  rom[38650] = 16'hffff;
  rom[38651] = 16'hffff;
  rom[38652] = 16'hffff;
  rom[38653] = 16'hffff;
  rom[38654] = 16'hffff;
  rom[38655] = 16'hffff;
  rom[38656] = 16'hffff;
  rom[38657] = 16'hffff;
  rom[38658] = 16'hffff;
  rom[38659] = 16'hffff;
  rom[38660] = 16'hffff;
  rom[38661] = 16'hffff;
  rom[38662] = 16'hffff;
  rom[38663] = 16'hffff;
  rom[38664] = 16'hffff;
  rom[38665] = 16'hffff;
  rom[38666] = 16'hffff;
  rom[38667] = 16'hffff;
  rom[38668] = 16'hffff;
  rom[38669] = 16'hffff;
  rom[38670] = 16'hffff;
  rom[38671] = 16'hffff;
  rom[38672] = 16'hffff;
  rom[38673] = 16'hffff;
  rom[38674] = 16'hffff;
  rom[38675] = 16'hffff;
  rom[38676] = 16'hffff;
  rom[38677] = 16'hffff;
  rom[38678] = 16'hff9d;
  rom[38679] = 16'h5263;
  rom[38680] = 16'hbd69;
  rom[38681] = 16'hf6eb;
  rom[38682] = 16'hff0a;
  rom[38683] = 16'hff2b;
  rom[38684] = 16'hf709;
  rom[38685] = 16'hf728;
  rom[38686] = 16'hff29;
  rom[38687] = 16'hff09;
  rom[38688] = 16'hff0b;
  rom[38689] = 16'hf729;
  rom[38690] = 16'hff49;
  rom[38691] = 16'hff28;
  rom[38692] = 16'hff29;
  rom[38693] = 16'hff28;
  rom[38694] = 16'hff29;
  rom[38695] = 16'hff28;
  rom[38696] = 16'hff29;
  rom[38697] = 16'hf72a;
  rom[38698] = 16'hff4c;
  rom[38699] = 16'hbd89;
  rom[38700] = 16'h5a21;
  rom[38701] = 16'hef19;
  rom[38702] = 16'hffff;
  rom[38703] = 16'hffff;
  rom[38704] = 16'hffff;
  rom[38705] = 16'hffff;
  rom[38706] = 16'hffff;
  rom[38707] = 16'hffff;
  rom[38708] = 16'hffff;
  rom[38709] = 16'hffff;
  rom[38710] = 16'hffff;
  rom[38711] = 16'hffff;
  rom[38712] = 16'hffff;
  rom[38713] = 16'hffff;
  rom[38714] = 16'hffff;
  rom[38715] = 16'hffff;
  rom[38716] = 16'hffff;
  rom[38717] = 16'hffff;
  rom[38718] = 16'hffff;
  rom[38719] = 16'hffff;
  rom[38720] = 16'hffff;
  rom[38721] = 16'hffff;
  rom[38722] = 16'hffff;
  rom[38723] = 16'hffff;
  rom[38724] = 16'hffff;
  rom[38725] = 16'hffff;
  rom[38726] = 16'hffff;
  rom[38727] = 16'hffff;
  rom[38728] = 16'hffff;
  rom[38729] = 16'hffff;
  rom[38730] = 16'hffff;
  rom[38731] = 16'hffff;
  rom[38732] = 16'hffff;
  rom[38733] = 16'hffff;
  rom[38734] = 16'hffff;
  rom[38735] = 16'hffff;
  rom[38736] = 16'hffff;
  rom[38737] = 16'hffff;
  rom[38738] = 16'hffff;
  rom[38739] = 16'hffff;
  rom[38740] = 16'hffff;
  rom[38741] = 16'hffff;
  rom[38742] = 16'hffff;
  rom[38743] = 16'hffff;
  rom[38744] = 16'hffff;
  rom[38745] = 16'hffff;
  rom[38746] = 16'hffff;
  rom[38747] = 16'hffff;
  rom[38748] = 16'hffff;
  rom[38749] = 16'hffff;
  rom[38750] = 16'hffff;
  rom[38751] = 16'hffff;
  rom[38752] = 16'hffff;
  rom[38753] = 16'hffff;
  rom[38754] = 16'hffff;
  rom[38755] = 16'hffff;
  rom[38756] = 16'hffff;
  rom[38757] = 16'hffff;
  rom[38758] = 16'hffff;
  rom[38759] = 16'hffff;
  rom[38760] = 16'hffff;
  rom[38761] = 16'hffff;
  rom[38762] = 16'hffff;
  rom[38763] = 16'hffff;
  rom[38764] = 16'hffff;
  rom[38765] = 16'hffff;
  rom[38766] = 16'hffff;
  rom[38767] = 16'hffff;
  rom[38768] = 16'hffff;
  rom[38769] = 16'hffff;
  rom[38770] = 16'hffff;
  rom[38771] = 16'hffff;
  rom[38772] = 16'hffff;
  rom[38773] = 16'hffff;
  rom[38774] = 16'hffff;
  rom[38775] = 16'hffff;
  rom[38776] = 16'hffff;
  rom[38777] = 16'hffff;
  rom[38778] = 16'hffff;
  rom[38779] = 16'hffff;
  rom[38780] = 16'hffff;
  rom[38781] = 16'hffff;
  rom[38782] = 16'hffff;
  rom[38783] = 16'hffff;
  rom[38784] = 16'hffff;
  rom[38785] = 16'hffff;
  rom[38786] = 16'hffff;
  rom[38787] = 16'hffff;
  rom[38788] = 16'hffff;
  rom[38789] = 16'hffff;
  rom[38790] = 16'hffff;
  rom[38791] = 16'hffff;
  rom[38792] = 16'hffff;
  rom[38793] = 16'hffff;
  rom[38794] = 16'hffff;
  rom[38795] = 16'hffff;
  rom[38796] = 16'hffff;
  rom[38797] = 16'hffff;
  rom[38798] = 16'hffff;
  rom[38799] = 16'hffff;
  rom[38800] = 16'hffff;
  rom[38801] = 16'hffff;
  rom[38802] = 16'hffff;
  rom[38803] = 16'hffff;
  rom[38804] = 16'hffff;
  rom[38805] = 16'hffff;
  rom[38806] = 16'hffff;
  rom[38807] = 16'hffff;
  rom[38808] = 16'hffff;
  rom[38809] = 16'hffff;
  rom[38810] = 16'hffff;
  rom[38811] = 16'hffff;
  rom[38812] = 16'hffff;
  rom[38813] = 16'hffff;
  rom[38814] = 16'hffff;
  rom[38815] = 16'hffff;
  rom[38816] = 16'hffff;
  rom[38817] = 16'hffff;
  rom[38818] = 16'hffff;
  rom[38819] = 16'hffff;
  rom[38820] = 16'hffff;
  rom[38821] = 16'hffff;
  rom[38822] = 16'hffff;
  rom[38823] = 16'hffff;
  rom[38824] = 16'hffff;
  rom[38825] = 16'hffff;
  rom[38826] = 16'hffff;
  rom[38827] = 16'hffff;
  rom[38828] = 16'hffff;
  rom[38829] = 16'hffff;
  rom[38830] = 16'hffff;
  rom[38831] = 16'hffff;
  rom[38832] = 16'hffff;
  rom[38833] = 16'hffff;
  rom[38834] = 16'hffff;
  rom[38835] = 16'hffff;
  rom[38836] = 16'hffff;
  rom[38837] = 16'hffff;
  rom[38838] = 16'hffff;
  rom[38839] = 16'hffff;
  rom[38840] = 16'hffff;
  rom[38841] = 16'hffff;
  rom[38842] = 16'hffff;
  rom[38843] = 16'hffff;
  rom[38844] = 16'hffff;
  rom[38845] = 16'hffff;
  rom[38846] = 16'hffff;
  rom[38847] = 16'hffff;
  rom[38848] = 16'hffff;
  rom[38849] = 16'hffff;
  rom[38850] = 16'hffff;
  rom[38851] = 16'hffff;
  rom[38852] = 16'hffff;
  rom[38853] = 16'hffff;
  rom[38854] = 16'hffff;
  rom[38855] = 16'hffff;
  rom[38856] = 16'hffff;
  rom[38857] = 16'hffff;
  rom[38858] = 16'hffff;
  rom[38859] = 16'hffff;
  rom[38860] = 16'hffff;
  rom[38861] = 16'hffff;
  rom[38862] = 16'hffff;
  rom[38863] = 16'hffff;
  rom[38864] = 16'hffff;
  rom[38865] = 16'hffff;
  rom[38866] = 16'hffff;
  rom[38867] = 16'hffff;
  rom[38868] = 16'hffff;
  rom[38869] = 16'hffff;
  rom[38870] = 16'hffff;
  rom[38871] = 16'hffff;
  rom[38872] = 16'hffff;
  rom[38873] = 16'hffff;
  rom[38874] = 16'hffff;
  rom[38875] = 16'hffff;
  rom[38876] = 16'hffdf;
  rom[38877] = 16'hffff;
  rom[38878] = 16'hffbe;
  rom[38879] = 16'hacf0;
  rom[38880] = 16'h7b65;
  rom[38881] = 16'hee8c;
  rom[38882] = 16'hff2b;
  rom[38883] = 16'hf72a;
  rom[38884] = 16'hf728;
  rom[38885] = 16'hf748;
  rom[38886] = 16'hf728;
  rom[38887] = 16'hff0a;
  rom[38888] = 16'hff0b;
  rom[38889] = 16'hff29;
  rom[38890] = 16'hf708;
  rom[38891] = 16'hff29;
  rom[38892] = 16'hff09;
  rom[38893] = 16'hff28;
  rom[38894] = 16'hf708;
  rom[38895] = 16'hff28;
  rom[38896] = 16'hf728;
  rom[38897] = 16'hff2a;
  rom[38898] = 16'heeea;
  rom[38899] = 16'hbd89;
  rom[38900] = 16'h5242;
  rom[38901] = 16'hf73a;
  rom[38902] = 16'hffff;
  rom[38903] = 16'hffff;
  rom[38904] = 16'hffff;
  rom[38905] = 16'hffff;
  rom[38906] = 16'hffff;
  rom[38907] = 16'hffff;
  rom[38908] = 16'hffff;
  rom[38909] = 16'hffff;
  rom[38910] = 16'hffff;
  rom[38911] = 16'hffff;
  rom[38912] = 16'hffff;
  rom[38913] = 16'hffff;
  rom[38914] = 16'hffff;
  rom[38915] = 16'hffff;
  rom[38916] = 16'hffff;
  rom[38917] = 16'hffff;
  rom[38918] = 16'hffff;
  rom[38919] = 16'hffff;
  rom[38920] = 16'hffff;
  rom[38921] = 16'hffff;
  rom[38922] = 16'hffff;
  rom[38923] = 16'hffff;
  rom[38924] = 16'hffff;
  rom[38925] = 16'hffff;
  rom[38926] = 16'hffff;
  rom[38927] = 16'hffff;
  rom[38928] = 16'hffff;
  rom[38929] = 16'hffff;
  rom[38930] = 16'hffff;
  rom[38931] = 16'hffff;
  rom[38932] = 16'hffff;
  rom[38933] = 16'hffff;
  rom[38934] = 16'hffff;
  rom[38935] = 16'hffff;
  rom[38936] = 16'hffff;
  rom[38937] = 16'hffff;
  rom[38938] = 16'hffff;
  rom[38939] = 16'hffff;
  rom[38940] = 16'hffff;
  rom[38941] = 16'hffff;
  rom[38942] = 16'hffff;
  rom[38943] = 16'hffff;
  rom[38944] = 16'hffff;
  rom[38945] = 16'hffff;
  rom[38946] = 16'hffff;
  rom[38947] = 16'hffff;
  rom[38948] = 16'hffff;
  rom[38949] = 16'hffff;
  rom[38950] = 16'hffff;
  rom[38951] = 16'hffff;
  rom[38952] = 16'hffff;
  rom[38953] = 16'hffff;
  rom[38954] = 16'hffff;
  rom[38955] = 16'hffff;
  rom[38956] = 16'hffff;
  rom[38957] = 16'hffff;
  rom[38958] = 16'hffff;
  rom[38959] = 16'hffff;
  rom[38960] = 16'hffff;
  rom[38961] = 16'hffff;
  rom[38962] = 16'hffff;
  rom[38963] = 16'hffff;
  rom[38964] = 16'hffff;
  rom[38965] = 16'hffff;
  rom[38966] = 16'hffff;
  rom[38967] = 16'hffff;
  rom[38968] = 16'hffff;
  rom[38969] = 16'hffff;
  rom[38970] = 16'hffff;
  rom[38971] = 16'hffff;
  rom[38972] = 16'hffff;
  rom[38973] = 16'hffff;
  rom[38974] = 16'hffff;
  rom[38975] = 16'hffff;
  rom[38976] = 16'hffff;
  rom[38977] = 16'hffff;
  rom[38978] = 16'hffff;
  rom[38979] = 16'hffff;
  rom[38980] = 16'hffff;
  rom[38981] = 16'hffff;
  rom[38982] = 16'hffff;
  rom[38983] = 16'hffff;
  rom[38984] = 16'hffff;
  rom[38985] = 16'hffff;
  rom[38986] = 16'hffff;
  rom[38987] = 16'hffff;
  rom[38988] = 16'hffff;
  rom[38989] = 16'hffff;
  rom[38990] = 16'hffff;
  rom[38991] = 16'hffff;
  rom[38992] = 16'hffff;
  rom[38993] = 16'hffff;
  rom[38994] = 16'hffff;
  rom[38995] = 16'hffff;
  rom[38996] = 16'hffff;
  rom[38997] = 16'hffff;
  rom[38998] = 16'hffff;
  rom[38999] = 16'hffff;
  rom[39000] = 16'hffff;
  rom[39001] = 16'hffff;
  rom[39002] = 16'hffff;
  rom[39003] = 16'hffff;
  rom[39004] = 16'hffff;
  rom[39005] = 16'hffff;
  rom[39006] = 16'hffff;
  rom[39007] = 16'hffff;
  rom[39008] = 16'hffff;
  rom[39009] = 16'hffff;
  rom[39010] = 16'hffff;
  rom[39011] = 16'hffff;
  rom[39012] = 16'hffff;
  rom[39013] = 16'hffff;
  rom[39014] = 16'hffff;
  rom[39015] = 16'hffff;
  rom[39016] = 16'hffff;
  rom[39017] = 16'hffff;
  rom[39018] = 16'hffff;
  rom[39019] = 16'hffff;
  rom[39020] = 16'hffff;
  rom[39021] = 16'hffff;
  rom[39022] = 16'hffff;
  rom[39023] = 16'hffff;
  rom[39024] = 16'hffff;
  rom[39025] = 16'hffff;
  rom[39026] = 16'hffff;
  rom[39027] = 16'hffff;
  rom[39028] = 16'hffff;
  rom[39029] = 16'hffff;
  rom[39030] = 16'hffff;
  rom[39031] = 16'hffff;
  rom[39032] = 16'hffff;
  rom[39033] = 16'hffff;
  rom[39034] = 16'hffff;
  rom[39035] = 16'hffff;
  rom[39036] = 16'hffff;
  rom[39037] = 16'hffff;
  rom[39038] = 16'hffff;
  rom[39039] = 16'hffff;
  rom[39040] = 16'hffff;
  rom[39041] = 16'hffff;
  rom[39042] = 16'hffff;
  rom[39043] = 16'hffff;
  rom[39044] = 16'hffff;
  rom[39045] = 16'hffff;
  rom[39046] = 16'hffff;
  rom[39047] = 16'hffff;
  rom[39048] = 16'hffff;
  rom[39049] = 16'hffff;
  rom[39050] = 16'hffff;
  rom[39051] = 16'hffff;
  rom[39052] = 16'hffff;
  rom[39053] = 16'hffff;
  rom[39054] = 16'hffff;
  rom[39055] = 16'hffff;
  rom[39056] = 16'hffff;
  rom[39057] = 16'hffff;
  rom[39058] = 16'hffff;
  rom[39059] = 16'hffff;
  rom[39060] = 16'hffff;
  rom[39061] = 16'hffff;
  rom[39062] = 16'hffff;
  rom[39063] = 16'hffff;
  rom[39064] = 16'hffff;
  rom[39065] = 16'hffff;
  rom[39066] = 16'hffff;
  rom[39067] = 16'hffff;
  rom[39068] = 16'hffff;
  rom[39069] = 16'hffff;
  rom[39070] = 16'hffff;
  rom[39071] = 16'hffff;
  rom[39072] = 16'hffff;
  rom[39073] = 16'hffff;
  rom[39074] = 16'hffff;
  rom[39075] = 16'hffdf;
  rom[39076] = 16'hffff;
  rom[39077] = 16'hffdf;
  rom[39078] = 16'hffff;
  rom[39079] = 16'he6fa;
  rom[39080] = 16'h7306;
  rom[39081] = 16'hc5ab;
  rom[39082] = 16'heeec;
  rom[39083] = 16'hf74a;
  rom[39084] = 16'hf769;
  rom[39085] = 16'hf747;
  rom[39086] = 16'hff2a;
  rom[39087] = 16'hff0a;
  rom[39088] = 16'hff2c;
  rom[39089] = 16'hf709;
  rom[39090] = 16'hff29;
  rom[39091] = 16'hff29;
  rom[39092] = 16'hff2a;
  rom[39093] = 16'hff28;
  rom[39094] = 16'hff28;
  rom[39095] = 16'hff27;
  rom[39096] = 16'hff49;
  rom[39097] = 16'hf70a;
  rom[39098] = 16'hff6e;
  rom[39099] = 16'had08;
  rom[39100] = 16'h6ae5;
  rom[39101] = 16'hef1a;
  rom[39102] = 16'hffff;
  rom[39103] = 16'hffff;
  rom[39104] = 16'hffff;
  rom[39105] = 16'hffff;
  rom[39106] = 16'hffff;
  rom[39107] = 16'hffff;
  rom[39108] = 16'hffff;
  rom[39109] = 16'hffff;
  rom[39110] = 16'hffff;
  rom[39111] = 16'hffff;
  rom[39112] = 16'hffff;
  rom[39113] = 16'hffff;
  rom[39114] = 16'hffff;
  rom[39115] = 16'hffff;
  rom[39116] = 16'hffff;
  rom[39117] = 16'hffff;
  rom[39118] = 16'hffff;
  rom[39119] = 16'hffff;
  rom[39120] = 16'hffff;
  rom[39121] = 16'hffff;
  rom[39122] = 16'hffff;
  rom[39123] = 16'hffff;
  rom[39124] = 16'hffff;
  rom[39125] = 16'hffff;
  rom[39126] = 16'hffff;
  rom[39127] = 16'hffff;
  rom[39128] = 16'hffff;
  rom[39129] = 16'hffff;
  rom[39130] = 16'hffff;
  rom[39131] = 16'hffff;
  rom[39132] = 16'hffff;
  rom[39133] = 16'hffff;
  rom[39134] = 16'hffff;
  rom[39135] = 16'hffff;
  rom[39136] = 16'hffff;
  rom[39137] = 16'hffff;
  rom[39138] = 16'hffff;
  rom[39139] = 16'hffff;
  rom[39140] = 16'hffff;
  rom[39141] = 16'hffff;
  rom[39142] = 16'hffff;
  rom[39143] = 16'hffff;
  rom[39144] = 16'hffff;
  rom[39145] = 16'hffff;
  rom[39146] = 16'hffff;
  rom[39147] = 16'hffff;
  rom[39148] = 16'hffff;
  rom[39149] = 16'hffff;
  rom[39150] = 16'hffff;
  rom[39151] = 16'hffff;
  rom[39152] = 16'hffff;
  rom[39153] = 16'hffff;
  rom[39154] = 16'hffff;
  rom[39155] = 16'hffff;
  rom[39156] = 16'hffff;
  rom[39157] = 16'hffff;
  rom[39158] = 16'hffff;
  rom[39159] = 16'hffff;
  rom[39160] = 16'hffff;
  rom[39161] = 16'hffff;
  rom[39162] = 16'hffff;
  rom[39163] = 16'hffff;
  rom[39164] = 16'hffff;
  rom[39165] = 16'hffff;
  rom[39166] = 16'hffff;
  rom[39167] = 16'hffff;
  rom[39168] = 16'hffff;
  rom[39169] = 16'hffff;
  rom[39170] = 16'hffff;
  rom[39171] = 16'hffff;
  rom[39172] = 16'hffff;
  rom[39173] = 16'hffff;
  rom[39174] = 16'hffff;
  rom[39175] = 16'hffff;
  rom[39176] = 16'hffff;
  rom[39177] = 16'hffff;
  rom[39178] = 16'hffff;
  rom[39179] = 16'hffff;
  rom[39180] = 16'hffff;
  rom[39181] = 16'hffff;
  rom[39182] = 16'hffff;
  rom[39183] = 16'hffff;
  rom[39184] = 16'hffff;
  rom[39185] = 16'hffff;
  rom[39186] = 16'hffff;
  rom[39187] = 16'hffff;
  rom[39188] = 16'hffff;
  rom[39189] = 16'hffff;
  rom[39190] = 16'hffff;
  rom[39191] = 16'hffff;
  rom[39192] = 16'hffff;
  rom[39193] = 16'hffff;
  rom[39194] = 16'hffff;
  rom[39195] = 16'hffff;
  rom[39196] = 16'hffff;
  rom[39197] = 16'hffff;
  rom[39198] = 16'hffff;
  rom[39199] = 16'hffff;
  rom[39200] = 16'hffff;
  rom[39201] = 16'hffff;
  rom[39202] = 16'hffff;
  rom[39203] = 16'hffff;
  rom[39204] = 16'hffff;
  rom[39205] = 16'hffff;
  rom[39206] = 16'hffff;
  rom[39207] = 16'hffff;
  rom[39208] = 16'hffff;
  rom[39209] = 16'hffff;
  rom[39210] = 16'hffff;
  rom[39211] = 16'hffff;
  rom[39212] = 16'hffff;
  rom[39213] = 16'hffff;
  rom[39214] = 16'hffff;
  rom[39215] = 16'hffff;
  rom[39216] = 16'hffff;
  rom[39217] = 16'hffff;
  rom[39218] = 16'hffff;
  rom[39219] = 16'hffff;
  rom[39220] = 16'hffff;
  rom[39221] = 16'hffff;
  rom[39222] = 16'hffff;
  rom[39223] = 16'hffff;
  rom[39224] = 16'hffff;
  rom[39225] = 16'hffff;
  rom[39226] = 16'hffff;
  rom[39227] = 16'hffff;
  rom[39228] = 16'hffff;
  rom[39229] = 16'hffff;
  rom[39230] = 16'hffff;
  rom[39231] = 16'hffff;
  rom[39232] = 16'hffff;
  rom[39233] = 16'hffff;
  rom[39234] = 16'hffff;
  rom[39235] = 16'hffff;
  rom[39236] = 16'hffff;
  rom[39237] = 16'hffff;
  rom[39238] = 16'hffff;
  rom[39239] = 16'hffff;
  rom[39240] = 16'hffff;
  rom[39241] = 16'hffff;
  rom[39242] = 16'hffff;
  rom[39243] = 16'hffff;
  rom[39244] = 16'hffff;
  rom[39245] = 16'hffff;
  rom[39246] = 16'hffff;
  rom[39247] = 16'hffff;
  rom[39248] = 16'hffff;
  rom[39249] = 16'hffff;
  rom[39250] = 16'hffff;
  rom[39251] = 16'hffff;
  rom[39252] = 16'hffff;
  rom[39253] = 16'hffff;
  rom[39254] = 16'hffff;
  rom[39255] = 16'hffff;
  rom[39256] = 16'hffff;
  rom[39257] = 16'hffff;
  rom[39258] = 16'hffff;
  rom[39259] = 16'hffff;
  rom[39260] = 16'hffff;
  rom[39261] = 16'hffff;
  rom[39262] = 16'hffff;
  rom[39263] = 16'hffff;
  rom[39264] = 16'hffff;
  rom[39265] = 16'hffff;
  rom[39266] = 16'hffff;
  rom[39267] = 16'hffff;
  rom[39268] = 16'hffff;
  rom[39269] = 16'hffff;
  rom[39270] = 16'hffff;
  rom[39271] = 16'hffff;
  rom[39272] = 16'hffff;
  rom[39273] = 16'hffff;
  rom[39274] = 16'hffff;
  rom[39275] = 16'hffff;
  rom[39276] = 16'hffff;
  rom[39277] = 16'hffff;
  rom[39278] = 16'hffff;
  rom[39279] = 16'hffdf;
  rom[39280] = 16'h9c6e;
  rom[39281] = 16'h6ac4;
  rom[39282] = 16'he68e;
  rom[39283] = 16'heecb;
  rom[39284] = 16'hf769;
  rom[39285] = 16'hf748;
  rom[39286] = 16'hff08;
  rom[39287] = 16'hff0b;
  rom[39288] = 16'hf6ea;
  rom[39289] = 16'hff29;
  rom[39290] = 16'hf708;
  rom[39291] = 16'hff29;
  rom[39292] = 16'hf709;
  rom[39293] = 16'hff28;
  rom[39294] = 16'hff27;
  rom[39295] = 16'hff28;
  rom[39296] = 16'hf729;
  rom[39297] = 16'hf72c;
  rom[39298] = 16'he6ac;
  rom[39299] = 16'ha4e9;
  rom[39300] = 16'h6307;
  rom[39301] = 16'hf75b;
  rom[39302] = 16'hffff;
  rom[39303] = 16'hffff;
  rom[39304] = 16'hffff;
  rom[39305] = 16'hffff;
  rom[39306] = 16'hffff;
  rom[39307] = 16'hffff;
  rom[39308] = 16'hffff;
  rom[39309] = 16'hffff;
  rom[39310] = 16'hffff;
  rom[39311] = 16'hffff;
  rom[39312] = 16'hffff;
  rom[39313] = 16'hffff;
  rom[39314] = 16'hffff;
  rom[39315] = 16'hffff;
  rom[39316] = 16'hffff;
  rom[39317] = 16'hffff;
  rom[39318] = 16'hffff;
  rom[39319] = 16'hffff;
  rom[39320] = 16'hffff;
  rom[39321] = 16'hffff;
  rom[39322] = 16'hffff;
  rom[39323] = 16'hffff;
  rom[39324] = 16'hffff;
  rom[39325] = 16'hffff;
  rom[39326] = 16'hffff;
  rom[39327] = 16'hffff;
  rom[39328] = 16'hffff;
  rom[39329] = 16'hffff;
  rom[39330] = 16'hffff;
  rom[39331] = 16'hffff;
  rom[39332] = 16'hffff;
  rom[39333] = 16'hffff;
  rom[39334] = 16'hffff;
  rom[39335] = 16'hffff;
  rom[39336] = 16'hffff;
  rom[39337] = 16'hffff;
  rom[39338] = 16'hffff;
  rom[39339] = 16'hffff;
  rom[39340] = 16'hffff;
  rom[39341] = 16'hffff;
  rom[39342] = 16'hffff;
  rom[39343] = 16'hffff;
  rom[39344] = 16'hffff;
  rom[39345] = 16'hffff;
  rom[39346] = 16'hffff;
  rom[39347] = 16'hffff;
  rom[39348] = 16'hffff;
  rom[39349] = 16'hffff;
  rom[39350] = 16'hffff;
  rom[39351] = 16'hffff;
  rom[39352] = 16'hffff;
  rom[39353] = 16'hffff;
  rom[39354] = 16'hffff;
  rom[39355] = 16'hffff;
  rom[39356] = 16'hffff;
  rom[39357] = 16'hffff;
  rom[39358] = 16'hffff;
  rom[39359] = 16'hffff;
  rom[39360] = 16'hffff;
  rom[39361] = 16'hffff;
  rom[39362] = 16'hffff;
  rom[39363] = 16'hffff;
  rom[39364] = 16'hffff;
  rom[39365] = 16'hffff;
  rom[39366] = 16'hffff;
  rom[39367] = 16'hffff;
  rom[39368] = 16'hffff;
  rom[39369] = 16'hffff;
  rom[39370] = 16'hffff;
  rom[39371] = 16'hffff;
  rom[39372] = 16'hffff;
  rom[39373] = 16'hffff;
  rom[39374] = 16'hffff;
  rom[39375] = 16'hffff;
  rom[39376] = 16'hffff;
  rom[39377] = 16'hffff;
  rom[39378] = 16'hffff;
  rom[39379] = 16'hffff;
  rom[39380] = 16'hffff;
  rom[39381] = 16'hffff;
  rom[39382] = 16'hffff;
  rom[39383] = 16'hffff;
  rom[39384] = 16'hffff;
  rom[39385] = 16'hffff;
  rom[39386] = 16'hffff;
  rom[39387] = 16'hffff;
  rom[39388] = 16'hffff;
  rom[39389] = 16'hffff;
  rom[39390] = 16'hffff;
  rom[39391] = 16'hffff;
  rom[39392] = 16'hffff;
  rom[39393] = 16'hffff;
  rom[39394] = 16'hffff;
  rom[39395] = 16'hffff;
  rom[39396] = 16'hffff;
  rom[39397] = 16'hffff;
  rom[39398] = 16'hffff;
  rom[39399] = 16'hffff;
  rom[39400] = 16'hffff;
  rom[39401] = 16'hffff;
  rom[39402] = 16'hffff;
  rom[39403] = 16'hffff;
  rom[39404] = 16'hffff;
  rom[39405] = 16'hffff;
  rom[39406] = 16'hffff;
  rom[39407] = 16'hffff;
  rom[39408] = 16'hffff;
  rom[39409] = 16'hffff;
  rom[39410] = 16'hffff;
  rom[39411] = 16'hffff;
  rom[39412] = 16'hffff;
  rom[39413] = 16'hffff;
  rom[39414] = 16'hffff;
  rom[39415] = 16'hffff;
  rom[39416] = 16'hffff;
  rom[39417] = 16'hffff;
  rom[39418] = 16'hffff;
  rom[39419] = 16'hffff;
  rom[39420] = 16'hffff;
  rom[39421] = 16'hffff;
  rom[39422] = 16'hffff;
  rom[39423] = 16'hffff;
  rom[39424] = 16'hffff;
  rom[39425] = 16'hffff;
  rom[39426] = 16'hffff;
  rom[39427] = 16'hffff;
  rom[39428] = 16'hffff;
  rom[39429] = 16'hffff;
  rom[39430] = 16'hffff;
  rom[39431] = 16'hffff;
  rom[39432] = 16'hffff;
  rom[39433] = 16'hffff;
  rom[39434] = 16'hffff;
  rom[39435] = 16'hffff;
  rom[39436] = 16'hffff;
  rom[39437] = 16'hffff;
  rom[39438] = 16'hffff;
  rom[39439] = 16'hffff;
  rom[39440] = 16'hffff;
  rom[39441] = 16'hffff;
  rom[39442] = 16'hffff;
  rom[39443] = 16'hffff;
  rom[39444] = 16'hffff;
  rom[39445] = 16'hffff;
  rom[39446] = 16'hffff;
  rom[39447] = 16'hffff;
  rom[39448] = 16'hffff;
  rom[39449] = 16'hffff;
  rom[39450] = 16'hffff;
  rom[39451] = 16'hffff;
  rom[39452] = 16'hffff;
  rom[39453] = 16'hffff;
  rom[39454] = 16'hffff;
  rom[39455] = 16'hffff;
  rom[39456] = 16'hffff;
  rom[39457] = 16'hffff;
  rom[39458] = 16'hffff;
  rom[39459] = 16'hffff;
  rom[39460] = 16'hffff;
  rom[39461] = 16'hffff;
  rom[39462] = 16'hffff;
  rom[39463] = 16'hffff;
  rom[39464] = 16'hffff;
  rom[39465] = 16'hffff;
  rom[39466] = 16'hffff;
  rom[39467] = 16'hffff;
  rom[39468] = 16'hffff;
  rom[39469] = 16'hffff;
  rom[39470] = 16'hffff;
  rom[39471] = 16'hffff;
  rom[39472] = 16'hffff;
  rom[39473] = 16'hffff;
  rom[39474] = 16'hffff;
  rom[39475] = 16'hffff;
  rom[39476] = 16'hffff;
  rom[39477] = 16'hffff;
  rom[39478] = 16'hffff;
  rom[39479] = 16'hffff;
  rom[39480] = 16'he6d9;
  rom[39481] = 16'h62a6;
  rom[39482] = 16'ha469;
  rom[39483] = 16'hff4f;
  rom[39484] = 16'hef0a;
  rom[39485] = 16'hf748;
  rom[39486] = 16'hff49;
  rom[39487] = 16'hff0a;
  rom[39488] = 16'hff0a;
  rom[39489] = 16'hff29;
  rom[39490] = 16'hff29;
  rom[39491] = 16'hff29;
  rom[39492] = 16'hff2a;
  rom[39493] = 16'hff28;
  rom[39494] = 16'hff28;
  rom[39495] = 16'hff28;
  rom[39496] = 16'hff2a;
  rom[39497] = 16'hf72d;
  rom[39498] = 16'he68e;
  rom[39499] = 16'h6b24;
  rom[39500] = 16'hbd93;
  rom[39501] = 16'hffde;
  rom[39502] = 16'hffff;
  rom[39503] = 16'hffff;
  rom[39504] = 16'hffff;
  rom[39505] = 16'hffff;
  rom[39506] = 16'hffff;
  rom[39507] = 16'hffff;
  rom[39508] = 16'hffff;
  rom[39509] = 16'hffff;
  rom[39510] = 16'hffff;
  rom[39511] = 16'hffff;
  rom[39512] = 16'hffff;
  rom[39513] = 16'hffff;
  rom[39514] = 16'hffff;
  rom[39515] = 16'hffff;
  rom[39516] = 16'hffff;
  rom[39517] = 16'hffff;
  rom[39518] = 16'hffff;
  rom[39519] = 16'hffff;
  rom[39520] = 16'hffff;
  rom[39521] = 16'hffff;
  rom[39522] = 16'hffff;
  rom[39523] = 16'hffff;
  rom[39524] = 16'hffff;
  rom[39525] = 16'hffff;
  rom[39526] = 16'hffff;
  rom[39527] = 16'hffff;
  rom[39528] = 16'hffff;
  rom[39529] = 16'hffff;
  rom[39530] = 16'hffff;
  rom[39531] = 16'hffff;
  rom[39532] = 16'hffff;
  rom[39533] = 16'hffff;
  rom[39534] = 16'hffff;
  rom[39535] = 16'hffff;
  rom[39536] = 16'hffff;
  rom[39537] = 16'hffff;
  rom[39538] = 16'hffff;
  rom[39539] = 16'hffff;
  rom[39540] = 16'hffff;
  rom[39541] = 16'hffff;
  rom[39542] = 16'hffff;
  rom[39543] = 16'hffff;
  rom[39544] = 16'hffff;
  rom[39545] = 16'hffff;
  rom[39546] = 16'hffff;
  rom[39547] = 16'hffff;
  rom[39548] = 16'hffff;
  rom[39549] = 16'hffff;
  rom[39550] = 16'hffff;
  rom[39551] = 16'hffff;
  rom[39552] = 16'hffff;
  rom[39553] = 16'hffff;
  rom[39554] = 16'hffff;
  rom[39555] = 16'hffff;
  rom[39556] = 16'hffff;
  rom[39557] = 16'hffff;
  rom[39558] = 16'hffff;
  rom[39559] = 16'hffff;
  rom[39560] = 16'hffff;
  rom[39561] = 16'hffff;
  rom[39562] = 16'hffff;
  rom[39563] = 16'hffff;
  rom[39564] = 16'hffff;
  rom[39565] = 16'hffff;
  rom[39566] = 16'hffff;
  rom[39567] = 16'hffff;
  rom[39568] = 16'hffff;
  rom[39569] = 16'hffff;
  rom[39570] = 16'hffff;
  rom[39571] = 16'hffff;
  rom[39572] = 16'hffff;
  rom[39573] = 16'hffff;
  rom[39574] = 16'hffff;
  rom[39575] = 16'hffff;
  rom[39576] = 16'hffff;
  rom[39577] = 16'hffff;
  rom[39578] = 16'hffff;
  rom[39579] = 16'hffff;
  rom[39580] = 16'hffff;
  rom[39581] = 16'hffff;
  rom[39582] = 16'hffff;
  rom[39583] = 16'hffff;
  rom[39584] = 16'hffff;
  rom[39585] = 16'hffff;
  rom[39586] = 16'hffff;
  rom[39587] = 16'hffff;
  rom[39588] = 16'hffff;
  rom[39589] = 16'hffff;
  rom[39590] = 16'hffff;
  rom[39591] = 16'hffff;
  rom[39592] = 16'hffff;
  rom[39593] = 16'hffff;
  rom[39594] = 16'hffff;
  rom[39595] = 16'hffff;
  rom[39596] = 16'hffff;
  rom[39597] = 16'hffff;
  rom[39598] = 16'hffff;
  rom[39599] = 16'hffff;
  rom[39600] = 16'hffff;
  rom[39601] = 16'hffff;
  rom[39602] = 16'hffff;
  rom[39603] = 16'hffff;
  rom[39604] = 16'hffff;
  rom[39605] = 16'hffff;
  rom[39606] = 16'hffff;
  rom[39607] = 16'hffff;
  rom[39608] = 16'hffff;
  rom[39609] = 16'hffff;
  rom[39610] = 16'hffff;
  rom[39611] = 16'hffff;
  rom[39612] = 16'hffff;
  rom[39613] = 16'hffff;
  rom[39614] = 16'hffff;
  rom[39615] = 16'hffff;
  rom[39616] = 16'hffff;
  rom[39617] = 16'hffff;
  rom[39618] = 16'hffff;
  rom[39619] = 16'hffff;
  rom[39620] = 16'hffff;
  rom[39621] = 16'hffff;
  rom[39622] = 16'hffff;
  rom[39623] = 16'hffff;
  rom[39624] = 16'hffff;
  rom[39625] = 16'hffff;
  rom[39626] = 16'hffff;
  rom[39627] = 16'hffff;
  rom[39628] = 16'hffff;
  rom[39629] = 16'hffff;
  rom[39630] = 16'hffff;
  rom[39631] = 16'hffff;
  rom[39632] = 16'hffff;
  rom[39633] = 16'hffff;
  rom[39634] = 16'hffff;
  rom[39635] = 16'hffff;
  rom[39636] = 16'hffff;
  rom[39637] = 16'hffff;
  rom[39638] = 16'hffff;
  rom[39639] = 16'hffff;
  rom[39640] = 16'hffff;
  rom[39641] = 16'hffff;
  rom[39642] = 16'hffff;
  rom[39643] = 16'hffff;
  rom[39644] = 16'hffff;
  rom[39645] = 16'hffff;
  rom[39646] = 16'hffff;
  rom[39647] = 16'hffff;
  rom[39648] = 16'hffff;
  rom[39649] = 16'hffff;
  rom[39650] = 16'hffff;
  rom[39651] = 16'hffff;
  rom[39652] = 16'hffff;
  rom[39653] = 16'hffff;
  rom[39654] = 16'hffff;
  rom[39655] = 16'hffff;
  rom[39656] = 16'hffff;
  rom[39657] = 16'hffff;
  rom[39658] = 16'hffff;
  rom[39659] = 16'hffff;
  rom[39660] = 16'hffff;
  rom[39661] = 16'hffff;
  rom[39662] = 16'hffff;
  rom[39663] = 16'hffff;
  rom[39664] = 16'hffff;
  rom[39665] = 16'hffff;
  rom[39666] = 16'hffff;
  rom[39667] = 16'hffff;
  rom[39668] = 16'hffff;
  rom[39669] = 16'hffff;
  rom[39670] = 16'hffff;
  rom[39671] = 16'hffff;
  rom[39672] = 16'hffff;
  rom[39673] = 16'hffff;
  rom[39674] = 16'hffff;
  rom[39675] = 16'hffff;
  rom[39676] = 16'hffdf;
  rom[39677] = 16'hffff;
  rom[39678] = 16'hffff;
  rom[39679] = 16'hffff;
  rom[39680] = 16'hfffe;
  rom[39681] = 16'hc573;
  rom[39682] = 16'h62a4;
  rom[39683] = 16'hcded;
  rom[39684] = 16'hef2b;
  rom[39685] = 16'hf749;
  rom[39686] = 16'hf729;
  rom[39687] = 16'hff09;
  rom[39688] = 16'hfee9;
  rom[39689] = 16'hff29;
  rom[39690] = 16'hf708;
  rom[39691] = 16'hff29;
  rom[39692] = 16'hff09;
  rom[39693] = 16'hff28;
  rom[39694] = 16'hf727;
  rom[39695] = 16'hff28;
  rom[39696] = 16'hff2b;
  rom[39697] = 16'heecd;
  rom[39698] = 16'ha4c9;
  rom[39699] = 16'h7326;
  rom[39700] = 16'hff7c;
  rom[39701] = 16'hffff;
  rom[39702] = 16'hffff;
  rom[39703] = 16'hffff;
  rom[39704] = 16'hffff;
  rom[39705] = 16'hffff;
  rom[39706] = 16'hffff;
  rom[39707] = 16'hffff;
  rom[39708] = 16'hffff;
  rom[39709] = 16'hffff;
  rom[39710] = 16'hffff;
  rom[39711] = 16'hffff;
  rom[39712] = 16'hffff;
  rom[39713] = 16'hffff;
  rom[39714] = 16'hffff;
  rom[39715] = 16'hffff;
  rom[39716] = 16'hffff;
  rom[39717] = 16'hffff;
  rom[39718] = 16'hffff;
  rom[39719] = 16'hffff;
  rom[39720] = 16'hffff;
  rom[39721] = 16'hffff;
  rom[39722] = 16'hffff;
  rom[39723] = 16'hffff;
  rom[39724] = 16'hffff;
  rom[39725] = 16'hffff;
  rom[39726] = 16'hffff;
  rom[39727] = 16'hffff;
  rom[39728] = 16'hffff;
  rom[39729] = 16'hffff;
  rom[39730] = 16'hffff;
  rom[39731] = 16'hffff;
  rom[39732] = 16'hffff;
  rom[39733] = 16'hffff;
  rom[39734] = 16'hffff;
  rom[39735] = 16'hffff;
  rom[39736] = 16'hffff;
  rom[39737] = 16'hffff;
  rom[39738] = 16'hffff;
  rom[39739] = 16'hffff;
  rom[39740] = 16'hffff;
  rom[39741] = 16'hffff;
  rom[39742] = 16'hffff;
  rom[39743] = 16'hffff;
  rom[39744] = 16'hffff;
  rom[39745] = 16'hffff;
  rom[39746] = 16'hffff;
  rom[39747] = 16'hffff;
  rom[39748] = 16'hffff;
  rom[39749] = 16'hffff;
  rom[39750] = 16'hffff;
  rom[39751] = 16'hffff;
  rom[39752] = 16'hffff;
  rom[39753] = 16'hffff;
  rom[39754] = 16'hffff;
  rom[39755] = 16'hffff;
  rom[39756] = 16'hffff;
  rom[39757] = 16'hffff;
  rom[39758] = 16'hffff;
  rom[39759] = 16'hffff;
  rom[39760] = 16'hffff;
  rom[39761] = 16'hffff;
  rom[39762] = 16'hffff;
  rom[39763] = 16'hffff;
  rom[39764] = 16'hffff;
  rom[39765] = 16'hffff;
  rom[39766] = 16'hffff;
  rom[39767] = 16'hffff;
  rom[39768] = 16'hffff;
  rom[39769] = 16'hffff;
  rom[39770] = 16'hffff;
  rom[39771] = 16'hffff;
  rom[39772] = 16'hffff;
  rom[39773] = 16'hffff;
  rom[39774] = 16'hffff;
  rom[39775] = 16'hffff;
  rom[39776] = 16'hffff;
  rom[39777] = 16'hffff;
  rom[39778] = 16'hffff;
  rom[39779] = 16'hffff;
  rom[39780] = 16'hffff;
  rom[39781] = 16'hffff;
  rom[39782] = 16'hffff;
  rom[39783] = 16'hffff;
  rom[39784] = 16'hffff;
  rom[39785] = 16'hffff;
  rom[39786] = 16'hffff;
  rom[39787] = 16'hffff;
  rom[39788] = 16'hffff;
  rom[39789] = 16'hffff;
  rom[39790] = 16'hffff;
  rom[39791] = 16'hffff;
  rom[39792] = 16'hffff;
  rom[39793] = 16'hffff;
  rom[39794] = 16'hffff;
  rom[39795] = 16'hffff;
  rom[39796] = 16'hffff;
  rom[39797] = 16'hffff;
  rom[39798] = 16'hffff;
  rom[39799] = 16'hffff;
  rom[39800] = 16'hffff;
  rom[39801] = 16'hffff;
  rom[39802] = 16'hffff;
  rom[39803] = 16'hffff;
  rom[39804] = 16'hffff;
  rom[39805] = 16'hffff;
  rom[39806] = 16'hffff;
  rom[39807] = 16'hffff;
  rom[39808] = 16'hffff;
  rom[39809] = 16'hffff;
  rom[39810] = 16'hffff;
  rom[39811] = 16'hffff;
  rom[39812] = 16'hffff;
  rom[39813] = 16'hffff;
  rom[39814] = 16'hffff;
  rom[39815] = 16'hffff;
  rom[39816] = 16'hffff;
  rom[39817] = 16'hffff;
  rom[39818] = 16'hffff;
  rom[39819] = 16'hffff;
  rom[39820] = 16'hffff;
  rom[39821] = 16'hffff;
  rom[39822] = 16'hffff;
  rom[39823] = 16'hffff;
  rom[39824] = 16'hffff;
  rom[39825] = 16'hffff;
  rom[39826] = 16'hffff;
  rom[39827] = 16'hffff;
  rom[39828] = 16'hffff;
  rom[39829] = 16'hffff;
  rom[39830] = 16'hffff;
  rom[39831] = 16'hffff;
  rom[39832] = 16'hffff;
  rom[39833] = 16'hffff;
  rom[39834] = 16'hffff;
  rom[39835] = 16'hffff;
  rom[39836] = 16'hffff;
  rom[39837] = 16'hffff;
  rom[39838] = 16'hffff;
  rom[39839] = 16'hffff;
  rom[39840] = 16'hffff;
  rom[39841] = 16'hffff;
  rom[39842] = 16'hffff;
  rom[39843] = 16'hffff;
  rom[39844] = 16'hffff;
  rom[39845] = 16'hffff;
  rom[39846] = 16'hffff;
  rom[39847] = 16'hffff;
  rom[39848] = 16'hffff;
  rom[39849] = 16'hffff;
  rom[39850] = 16'hffff;
  rom[39851] = 16'hffff;
  rom[39852] = 16'hffff;
  rom[39853] = 16'hffff;
  rom[39854] = 16'hffff;
  rom[39855] = 16'hffff;
  rom[39856] = 16'hffff;
  rom[39857] = 16'hffff;
  rom[39858] = 16'hffff;
  rom[39859] = 16'hffff;
  rom[39860] = 16'hffff;
  rom[39861] = 16'hffff;
  rom[39862] = 16'hffff;
  rom[39863] = 16'hffff;
  rom[39864] = 16'hffff;
  rom[39865] = 16'hffff;
  rom[39866] = 16'hffff;
  rom[39867] = 16'hffff;
  rom[39868] = 16'hffff;
  rom[39869] = 16'hffff;
  rom[39870] = 16'hffff;
  rom[39871] = 16'hffff;
  rom[39872] = 16'hffff;
  rom[39873] = 16'hffff;
  rom[39874] = 16'hffff;
  rom[39875] = 16'hffff;
  rom[39876] = 16'hffff;
  rom[39877] = 16'hffff;
  rom[39878] = 16'hffff;
  rom[39879] = 16'hfffe;
  rom[39880] = 16'hffff;
  rom[39881] = 16'hffbd;
  rom[39882] = 16'ha46d;
  rom[39883] = 16'h7324;
  rom[39884] = 16'hd64a;
  rom[39885] = 16'hef2a;
  rom[39886] = 16'hf729;
  rom[39887] = 16'hf708;
  rom[39888] = 16'hff0a;
  rom[39889] = 16'hff29;
  rom[39890] = 16'hff29;
  rom[39891] = 16'hff28;
  rom[39892] = 16'hff2a;
  rom[39893] = 16'hff28;
  rom[39894] = 16'hff48;
  rom[39895] = 16'hff49;
  rom[39896] = 16'hf6ec;
  rom[39897] = 16'hbd49;
  rom[39898] = 16'h6ac3;
  rom[39899] = 16'hbd71;
  rom[39900] = 16'hffff;
  rom[39901] = 16'hffdf;
  rom[39902] = 16'hffff;
  rom[39903] = 16'hffff;
  rom[39904] = 16'hffff;
  rom[39905] = 16'hffff;
  rom[39906] = 16'hffff;
  rom[39907] = 16'hffff;
  rom[39908] = 16'hffff;
  rom[39909] = 16'hffff;
  rom[39910] = 16'hffff;
  rom[39911] = 16'hffff;
  rom[39912] = 16'hffff;
  rom[39913] = 16'hffff;
  rom[39914] = 16'hffff;
  rom[39915] = 16'hffff;
  rom[39916] = 16'hffff;
  rom[39917] = 16'hffff;
  rom[39918] = 16'hffff;
  rom[39919] = 16'hffff;
  rom[39920] = 16'hffff;
  rom[39921] = 16'hffff;
  rom[39922] = 16'hffff;
  rom[39923] = 16'hffff;
  rom[39924] = 16'hffff;
  rom[39925] = 16'hffff;
  rom[39926] = 16'hffff;
  rom[39927] = 16'hffff;
  rom[39928] = 16'hffff;
  rom[39929] = 16'hffff;
  rom[39930] = 16'hffff;
  rom[39931] = 16'hffff;
  rom[39932] = 16'hffff;
  rom[39933] = 16'hffff;
  rom[39934] = 16'hffff;
  rom[39935] = 16'hffff;
  rom[39936] = 16'hffff;
  rom[39937] = 16'hffff;
  rom[39938] = 16'hffff;
  rom[39939] = 16'hffff;
  rom[39940] = 16'hffff;
  rom[39941] = 16'hffff;
  rom[39942] = 16'hffff;
  rom[39943] = 16'hffff;
  rom[39944] = 16'hffff;
  rom[39945] = 16'hffff;
  rom[39946] = 16'hffff;
  rom[39947] = 16'hffff;
  rom[39948] = 16'hffff;
  rom[39949] = 16'hffff;
  rom[39950] = 16'hffff;
  rom[39951] = 16'hffff;
  rom[39952] = 16'hffff;
  rom[39953] = 16'hffff;
  rom[39954] = 16'hffff;
  rom[39955] = 16'hffff;
  rom[39956] = 16'hffff;
  rom[39957] = 16'hffff;
  rom[39958] = 16'hffff;
  rom[39959] = 16'hffff;
  rom[39960] = 16'hffff;
  rom[39961] = 16'hffff;
  rom[39962] = 16'hffff;
  rom[39963] = 16'hffff;
  rom[39964] = 16'hffff;
  rom[39965] = 16'hffff;
  rom[39966] = 16'hffff;
  rom[39967] = 16'hffff;
  rom[39968] = 16'hffff;
  rom[39969] = 16'hffff;
  rom[39970] = 16'hffff;
  rom[39971] = 16'hffff;
  rom[39972] = 16'hffff;
  rom[39973] = 16'hffff;
  rom[39974] = 16'hffff;
  rom[39975] = 16'hffff;
  rom[39976] = 16'hffff;
  rom[39977] = 16'hffff;
  rom[39978] = 16'hffff;
  rom[39979] = 16'hffff;
  rom[39980] = 16'hffff;
  rom[39981] = 16'hffff;
  rom[39982] = 16'hffff;
  rom[39983] = 16'hffff;
  rom[39984] = 16'hffff;
  rom[39985] = 16'hffff;
  rom[39986] = 16'hffff;
  rom[39987] = 16'hffff;
  rom[39988] = 16'hffff;
  rom[39989] = 16'hffff;
  rom[39990] = 16'hffff;
  rom[39991] = 16'hffff;
  rom[39992] = 16'hffff;
  rom[39993] = 16'hffff;
  rom[39994] = 16'hffff;
  rom[39995] = 16'hffff;
  rom[39996] = 16'hffff;
  rom[39997] = 16'hffff;
  rom[39998] = 16'hffff;
  rom[39999] = 16'hffff;
end

always @ (posedge clk)
begin
  dout <= rom[addr];
end

endmodule