//===================================================================================
//Author    : TRZ
//Data      : 2021/08/16
//Funcation : IO 滤波
//filter time = FILTER_CNT * (1/filter_clk) 
//===================================================================================

`timescale 1ns / 1ps

module	cb_filter_app #(
    parameter     OPT_NUM      =   40  ,
    parameter     FILTER_CNT   =   8   
)
(
//-----------------------------------------------------------------------------------
// Filter & System Clock & Reset
//-----------------------------------------------------------------------------------
    input                               filter_clk                  , 
    input                               sys_clk                     ,
    input                               rst_n                       ,  
//-----------------------------------------------------------------------------------
// Orign IO Photoelectric Signal input
//-----------------------------------------------------------------------------------
	input     [OPT_NUM - 1 : 0]         orign_opt_i                 , 
//-----------------------------------------------------------------------------------
// IO Photoelectric Signal output After filter
//-----------------------------------------------------------------------------------
	output    [OPT_NUM - 1 : 0]         filter_opt_o
); 
//=================================================================================//
// -----------------------------------Instance Area------------------------------- //
//=================================================================================//  

genvar		bit_num;
generate  
	for(bit_num = 0 ; bit_num < OPT_NUM ; bit_num = bit_num + 1)
        begin : IO_FILTER_APP 
            cb_io_filter # (
                .FILTER_CNT             (  FILTER_CNT             )  
            )
            U_cb_io_filter
            (
            //-----------------------------------------------------------------------------------
            // Filter & System Clock & Reset
            //-----------------------------------------------------------------------------------
                .filter_clk             (  filter_clk             ), 
                .sys_clk                (  sys_clk                ),
                .rst_n                  (  rst_n                  ),  
            //-----------------------------------------------------------------------------------
            // Orign IO Photoelectric Signal input
            //-----------------------------------------------------------------------------------
            	.orign_opt_i            (  orign_opt_i[bit_num]   ), 
            //-----------------------------------------------------------------------------------
            // IO Photoelectric Signal output After filter
            //-----------------------------------------------------------------------------------
            	.filter_opt_o           (  filter_opt_o[bit_num]  )
            ); 
		end 
endgenerate
  
	
endmodule 



